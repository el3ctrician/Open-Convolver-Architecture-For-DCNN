`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mJ+PLYjKLUXjMwYVEVUe0bjwKU4L557171yjEjJtGS7XYhYuTZ2EhxyPWOHTtB6rbJ7dNTpa4+GE
wBtjk1Yb2g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
KhNdPJEFiKsVcA3vhRwZ9mjxzSg0HP3McYNBsHeYxhzKDeIbU0QGJU/JsE9IK78cwUVGGyv7nosv
ShgEKqDGjEHTs5bChGs9DwyTOj91l50JWJYfJ0B+1z22kPchk4Fqpe/dA9NdiloMAYWh/G80o2l4
8J0b+l7MrhDRQwCLjUg=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
E/IWYvoiGjNzlk34mDFPjIvEGfsCMF5+MilbaIgK2K3aWG+Moimutsp4HT8zVy6YwSudB1axFp7L
Isza5I7Bq99mEc2S2PAqnH/GZlYJ57DmrrVV2SYLXCkWqUe9qyaX1CxVXQWNFS0VwSsIuT9qGQ5y
xKWC24LxF0GymDWhzPo=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QS2h/dgW5k9f+uPAGJgxFy52DUOQxnQ0E/v373wAdvAbJmE5aDq+hCiQpKjIy4GPR18nf0BhvZks
RspM6uNQT4RbJ0TuXkCg9Lpa0+6DHVRStYYifhXoayvXLRda/xPDCdRoWjyVDYwy31/VtVUUd4sk
WporoUtt67H4PtSQmJtPZpeIUrGdC+kxUF0hCSTPP0g74SGWqjJO6MYy2GpV1LkKC99zUdygglNt
NaN9lwF+nKe4Fg0FvdqhGv6N3nGeI1MJK6txjmhg954ucmXziIj4uwERSPXebVI8b/ZABz/VEbS9
VxBY/edTEMmjFBPAAyi4+nMCIBico/hk9209kA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pycQ2fLSVY13WgerGDIXIscwMlm8GzUI80lStjmrI+BFUJvWAeXjSGUMHboPoeLKC4wublBqYtsx
gt0DMJlDYdpjuptV0As8xM9hETwEA3wJtQZRmsnqGPE9m9JRCIQRD+xAicjW/zhztX16wJUIHtWx
l2WVqFeSzjUtrU/RogUILCxN0UcvYY8FdlRpjEF9WwNnZpz1vaFyrA2vYbE/Hb9Ir41wGK+zTWJs
gWEP3XuO3BPXTg4RaVK1UNC2cI/P8ovP1+2Ad8N5Sz/+dX+n/IZ0Q0TOE6fBmh8ZcbmwCxclw0jG
BQhscdUhX/wWXCxVGWwQX/CRuo+hYOuae1iNQg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mAQF9E53i8C7OIv2LDuX8SwOm8wguKByZfIGIplx/BUXP38mOp3CAXU0i43ZSjzf9p5bNnYAdA9T
SVTvziFLfJqU2HwQw4kLAXCTqpx/Kc5kV2cMGlzTB0UKNnSnjZPWTIE2pcMOfN+GXN4XUZ+/sHtE
e+UuO9YRuFV1zYpwtLtHM7EokzmoZDakqLb0EVzJMYXit7Kx9S8d3AwEoC5UGon7KtaLY9OSTPuo
EjbktSML1hmkbUGLhPFpp38+uxx8nTBWs6GJuTksSZf3lOWi9N+mWAvgw3PPhyPT/3ERw30zvMHz
TtsPw5PGrfcFsOmvqIBfVP/KSHUFfNnS9SyhOA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 261312)
`protect data_block
C7k/tG/ONC/2vI3YDtVI9fIUOZ2nDdVjDCTVJ4EnzGcjeY+ocM4zWh1DqEDnOu98kPulT1+dQJxN
fiPodHgiJgANI7bdY17a3gz0eRHXQlWUoYH5lVZyBB6ESClH3QezhN7R1f/XxvDxNw640l5HlcS/
0okKQBrRomfXREj1KCe9/KBdgwxcdAH1VveCM7wc1KEUbUUSWh91/9ZXCn/FV9IVguUA3D1HIkdw
CLorKhhIjbKyOdZitYY2wsRiv4q1cgRSala8I62h7E7o5Kbvn2Xu2aeNIzM4DDRfIlY703quix19
2A1uJCn3B1tiVpGcIYTFKwztgzWhd5s89B2/H8v4m5K8IaXEMpkW5EA4jVnCUPc0IHlZelcTJOhc
vCDWzQxpQVYHNYWX1wAHbGlsP9caOu8nwUEEUmI51g+lugrO1JcluBFm2smHRFEr9z+wj7zRiqsh
3o6/AkjKCOymNSrF76uQbDDGLxpBrcFDCtqTsQIn7V7tFEi4M3qTWflBvy+aF8Th9rTWsXIcP5SD
cd0CaijmZJ3GiDo4lCClmGRGH837H+lcfYolIBzSBJGUEgFiuynzFfwQh+0rlP5/FMlj+6bOB5Un
2RGMeORHP2DeVDYdQBg4wLRfJHWEPAlFzpaL/7zBLIuOLryFJVWJuBy0EzNO+XpflLvS9xSj8/YJ
XJAzh6536O/WxtX+9JAd9Ko6SMfvTdmJ54oja5IC/VorHDEeZdwBHFSv/LTl3gOnM0f/ZGt59jNo
hc833uFdKSfG8LJ4LAaoJPQwt02UmckGsWmEJmBnmWgdQkuOQHvMjx1o06jfurFuXtfdRrsaXJ9O
J7IehhTTmje4aTdVzVF6+Q2qszt4KHR2U4O5x5yHUC01cM/A/xWDJA34QBoUfMF5CvG3SgvrVi5s
KaJTVA43aTdJT5aPtvKAHelz3WUMEl3E8gJ9/3rBI50NSZNxuE14FAfDQZy8HyPOX+Yr8MALE23V
fk0UpdifitjTirMswEiFuXkrzoGTiCZP0cmBFmcKMBAR5le3pkNIpW1G416/2JimSDq4GnFrr7zW
wtHpHzQycikzg0fQTBjd0rsgEVd7aUhTTnxlqbyyZ+f5wWGYyJyNiGagw8+nJyZyliednl+IiIa4
my8Dfcx6f46en4iXdSi5Dt9BrdrSDsxC0jO9fzYv+HvRzESXFweGQQwaoGr+BtGaGkzoCAZ97xNQ
ABWjUuTZCpPrs2sPgCxsVEAXnphgIDsFfpg158g1nRsNZ7prCuphdgortG7f89ppwPkaP1Izh7oq
AylP6+dHLO4om80BqXFZrFMosbVhtrpdaHoESmpikHQpnxRW/0os2a9HF7vGaJUU//J/pJBiWn2P
+eArM51rY4HgEDJ3oD1smC8/7cXdG9ZMk0dKPK+P8SYBIY3cXqiMYwibONz1rYXiytfOQyN1cXTc
0Eir9W9YQyBZ0F/haAag2jIDVdLjZUuVl3J8dsJ5dbb9eYW/HAnLnEQK0ziIFW95cbbQWLBznZBj
MxQQjarTCEvlPqjGAV9miZ7hjq38/0E8+rWHAxkrDH2dsPbGIj+uvvztQwG2QwLv1Hrfd296Zzyo
gU6blkZS3wMdPvX8C5C2lc6Xg48feFZ3sZcrR0swhwKFsSCJ91DIqJGNbTmm4HRnCQBouPsLwN4p
1LEcurelyDHm2Yc/ZvlAjinFgc2v9zkfpddB0qI68FYqoJe5m5XPr9nrhngyea2dwZXH3QhUKHV2
ilKKcSvv/8GlVDdvabtgNpW0QrxSUPGlGy4S888uwMFO+gSwd+nyzdUTd9sgmqJG4WnNlbl4gkho
yxbuepxH2naO5Vd5+sPu3yHx8qxWWVKTV8BkDfIIfHhszfxMczZDM5kyD44lEARE4zAxmk/amQlH
U3j6muJ9QBrs/SUO7dEAeMUE/4ZXQP9zJhd+OIbJvgIBAb/26Olium6N2CtL9UZEvM5nxhjsB3Sl
schId/datpC7Z4vJHb0sy7DARsCjTWxBB0Qt6gQstXoKnthDdMp867ykMmZNpYtsoFkWwQLnS0mA
2B6HsFK9boXzUqz4Dmgf45XsNyLh+Cvrj8mW0ns1tbohSrcMmiDkd4A3cgEv9jyCIrqljTCYx91r
HaHBEDssVoqU/2PTh6Mpt5vQzHkrSs4oTuzDfpvtXYlFdCyZxkB+N5hNjvZdmnkeSXkKh5ElZi9w
NqlWZv5PQuRybGirwEWui7d7JhsKJPNNlAXe+Zm4h99efObdK6BsNsLNwD8daCaERkgY+6PeUVqU
39QguBaPpMnp6zjeuNBalUo/5vnBVSOUiAXoA/P1rUM9J7aGNS34GpYRXjJqFAg6rD4o4QJXpY2a
iAHbNZBw7ujEULHX5zyTVz/3rn8Z/EE6zlfGw3tcTH/rnTAcXk2Dkv4rbATi71JPp6E7MK/LnSxn
q+y7Sy0Rk2m68GK8WOeDubBE32vmPVQZEgq287KfLMQQbeTnwrFakPmxYeqkJ7uoOEvCPrf1iU4t
HkoB3CYAJuvT7RaXegIFxY6Z/hAsgLCW8WFZ1woaE6aomPAiXx5gIPLLINW014FyytF4YW05JtsL
XpZmhH/0pV4mtbHPM+LBICxdCD0NCVsRhQhclrz2yikRILYNBDLRpEhhSsq1ZdJjZkZc5S4DxeQS
4GwPnSCeOKG0xHTkE7sAzi6nnGBRtfua//ZdvndzMHvL92E8/iI4qhY6lCr45bBAkh2kCcxLfIbC
4AhLQJILmfeEil2/MFTvmsmU+7b0FALvgZkD640no6r3SQcssfFnTCx2cIcjh51F3tdPaRRzPk9y
ZsflsqIM5ejmQJKrmaQpkceDgkCYboqPyTpFM2lyhinoJk4w7RCjKZkZJdh1s4lem40+ZbrpSpjf
kX90z3jsdZZh/Nq9na4KQ1xsNwb3mjS1Vel6yiM9FU3P6qb5mMh434ezcxyRCQH0/RKTTAEyXRWx
1DUbnX38/VEU3RxvBPjlAo6TzbXZ4eaDzm86p4CSBQbhty237IEqut+Ck8yzNNRXlm5eYRlCyTFE
zLF4dskI87p86jod7qGYnu14QVrtmqEH61Ew9GGBzhvfIYKWs9wHMLx4EqTb3VPsn8ppES66U4K7
zc+j2jmKtzKM1egwUrJrQGdBFHBKBEdeCRjcyWaWycVHW9C5gf4CSAi8hj+rCDuWlXN8mqoZBf3p
Lu8+oiWwmQYeJhHmHXEkq/0GnBoKhXp3+w5z4blZmC2CeK3SysKoL5jKHj2Y1EuSUbRi3+U4jv7e
zD92bXq3XkkOJIdwzaK6PCP/cQDXWXu6rikzcvaWdh11IJuV7SKRQJjsSbEoFqpyUL9bBhobcEM2
wWiuwJr6x6NsGm/jB3p4va8m+5nVLz5LDDygyPOyiuqB/fym08fjOKtI7xMoRc94XhifKwbsjRJa
No22XXcMWhL1VMgVbxmWEsEEiuC8sZx0p1gDX4kEHEeI19fZLOF0aER/VWrUAfOa0SiISRJpPp7p
gsdle539Kp1+JiMR9Uv1XstikVYYlJnKH4rJhesaoAiZkGtx7BXTLAR/cLSF/XeuoBO5nx8aHEqV
2kg5HLWIxS/44MKWYSys2ElEI+swqVN5KtcFo7e8fX6WqjfjHI/Ee7Gl8ZqDKPKsxhWCkx5tm9r3
2QQ8qomtsVeyojy47pcfYhXjIVD6F3xTrB7YQrRI3ZpVasiymzd72E1wGlrzCamEiZuDLff9hLt/
WWB07GYcorfzxOzD5XyDwsQrQeZ/MGtCyHGfym5MBnnN8Gw9lV4KlITetubR8zf9qhsLIVpRhe/7
mkVHPk0Z2PabSKVMLLnw7St/uhTSWM8GulIru8BncNhK3bNoEzzZV0Obev517Yzacrk6nydu5BSs
QzqPCKCG3WWaH3ROTPG0CxjE1mcaCmeGdSkLMt4v44gwwJ7rrA0I4VajPk49Tr0VG25d5IiFa8Js
HKZWE8CMXqR2ycz6AdYT4XikDvxT7yDF3DbxybjA8abfUnUWBkHMQxZoUQKSXvq5+ql8iW0EcWUM
rW32ugLtgrw0+fAwngA989spwpDSiy02WnuRF1CdvIQKNcIEx2Wy4G/t3CZ7BBkj9gxYug2FVBmu
O87MWeJ9abe4v61BLxjcUxfDE6D+nB3QwPzV9qbmoXU4/aqFcgDHP6Rhb9ENe1YxfRTcVJosMKQo
zHbgKdYgUV1FxH5ZSUm3Jm14NQIl5K/Gs9URkXIOrVyyaf562CN5+pUq/CzEiQ5yyJWdPjTA3jpv
R7bZEDd46k3teMKWpYoKWfAR9FpnHmFMPezHqVJOodMNVyiOpBXQeYckLpnHN4fzfmTmQUqXkrs8
FQscwh7Fg13jJA1FpZfK9oCVqFuJJfXF0dnTYwKu46tPQJ98EtmGJo+pNyDMv1qeOv2MfoDtJrAh
xY98GPhg48mUjJ2TvnUQvWmjWakvgN74e1E0S1lCbeFCKib9RNd+mYWqj8nQY0QH+0VqEatRHTIn
jzaAvS5U9j1LzY6FXlUWXd5mXJ2pJS8ZS/+nXYZfqiQRGvNoel11b7lo3FNHvJ/L1KgkyM7e59Rz
gV9V5U/6bBoOwOfMjJjStX023hLk3m6zycKhV4D+46uQkPAE9X+gY6wFFbGLsmv2v5FNVflyjDf5
8gpFja9t/wnRP+kcYGkOx+zqTMZCNOwjbM8X8mM4iAhIfiuk0s/J7bqAOeqmKvTdjJBK9/8J85WB
3XMN3UBA5Ygu4JYEkwZwaCQd5WmE57UvpgaatPo0UWnOLmYqfsOfJbzsdUfowLZDkfIWvPsVmxcZ
fA1s9gxghC6LmLGZJ1Icg7EJuVum36KxBMXaOAyizpk+i0Xt2kdylmRhv+7myKEEER+wx+OC5oZv
VUlFAADKZk2hcb809UYzTbwr4CytObF2I3C6yi3UqpFS/y+9/UCAzAYkjSd0sc06+to4YUougNqN
NOdQsyGyAkPkKSEzLPocizKxAwr/luWM4olBRaaeqN+6umfGk/nflrjHHJtT3piXXfc1NDKz2Pyu
JrDr2lsVP+cgXKinO72FNqVsque7lXJdYv2xitCOvxxAVzMravi/b2llYGjqwy5UhUf/u6jL5JTE
jrvfLDKFBT5wNCnaIk1Vr5c26QWZ7C+UJafx0Z18tc7D9MrFucKh8btuHJt038/CQyPow6Dj9wjj
ASo3QG5EvN2TBbeuKzimm+jNfLMJd3orVEZx09C16+as2VIDaBo9/tLimc//RmGe7DElP+oBHiUh
bTqvIE3++eMfk6l7AEfWavEH/KeXjYylVFVFrnAJoenHqrtwms7K6d1q44itux/xZXv6Bb2YVArK
PLIjJJ52+wtmV0pGFBd7YQBh92dktz9KBuiDcRkJKOsnrD4BoygTGI0aMhzHWzJKF7uDBYnFoY+M
ixemw4YoP9v2DZCyfO77gvRU5kQluPkAqOP6E0UCjPVcoXV+AZ4r0qjh7mexxA5LcLW717tY3UAt
3rjwrQUydOhP6sM7chs+0aJ0zxZknVKbg/zg6JzZ9LtYXWBhSDkhSVPF2u6IRGuwgzLnzNOtTcsU
NYND72uq6l0z9U2FcVv+vi3KCspMTNqBtEOAt+XHQ5/WUju2v3/QPPuKVzO8iAuabK3GPQNywE3+
yxsbp0NHyOYjsB0uKVlyH3f1E2KXsqwv4q7vsVqwI3e0c6SltVFFrwNgNRrbPpRHP8+RwEQmxbz4
r7dUeqvy5tcK0UFqVVrlLQO5ILhHVsktY7TcbdptzkrkknnZAghQdDfKc10UGY4YqWMtF5MK+In1
/cRQt/kYkIPFkXS4ixKbPcsB+LaFYmM9uk31Qj67l2ENiiJZaWHvyMk29690JxZpDJzZhE5zZuel
P4Zi7iD4tmRnt7ra3XTfeqcjwpoFCBzw8SVYkPX7wicDdvIKSBTfzMjXCRZO0N2jWIALZI5M0WZr
JXUUFiWDxHgVWPJMw1bCZD29wCk5P6nlT9Wf8e+kw2levcph2RLmNdZmEUdsdL9EAoS4rSaveM9P
cliBD3rQnFruOd9eFSA/XbkBEiEc9x6UmJ7bcJvTsMeGea6DsVkj0bbQphcXh/9ItVMEMNsUQN/Y
+/qUnbENu1Bb0MMNzrRlgepJ9ovsbDPHaBKFLN042sa/pteK/SRu7MYw7iDN+uJBR6BK+9bAXNRm
X9STOa7TgcqzxOU+UDUBQj6vXa4jpa6YzxVLybt3v0yGZSsGlyETRHmILllIBBbvWUuW3GcUbV1s
EiPsaPy9i3Dn77ha94wGphEAW1ix0Vg0AL7DPrneH/6awjHxmD5RRiPKFbctXfpXqX5PHg+lD8eX
gbnWKOAEsQMq2q4u+SyrHk+JeEyd5VcheY/Jz/TMilUmdWXKY51Ab7d6um0ndfLKFOORDJHMXGAW
hI3j+JColozZGl1ETQzLHozOT18FGM5cUPWSKzkE8UPeBsOhz89+Ba2pN+m13Z3Wu6HcmnAMWcff
Sd9t/pljYIjgwYjMw5XQMyHhPmP6dRBu8KgJIPbr5VSn/5ATlD0qh9P2z1MOwwk3qrHZKxEl5l2g
tj2btmOLooVCZC2CEjsmR+LcgF+tszHweyZ0DGrtSbd2iXYy51r4tRjB/389xNYnbcBwmkuvZPRL
HwHem5y4Ov9T+MJcLLHh/8d/kpSS0Lv/8LR6AkxLO00a7KIZsVQIIDJlDQuTSjfvcpL+zDCySg2I
gkHIN3wW1D9Lk39eDmasiQs1eXF0CwKHQzGerodzYRQTdCcr6uArUSkXZIRI/ZEQW3ncZscHWnDt
dZPivhxX3/18gcSAhI+KYNhlBkmlWiKFwJs1UxH6pUguJ609Ckq1h/1eFLD1z8wXJQeZjs8ARHvl
gnwLnxCjmb/rU88OOch0K55p3hEVXjrGgIBDqffgEEYhN9qUbieIUOkcsih6cJHzK0Opx65lRr2T
ktOgEo4WCFVvSuZ/zSe4WZvPsll9uQDogzgsr2+gG8ogqFkqMdgar44eQUOsV5Ew4ZYVkeZKnheV
w0+Rmc3KmzwRnQpWtELv2BnWcwTP74rWdlskNNJC9pZ2VxzywNVYKIhyc/7xxgd4l6uqC+FT4cO+
Xg/w5dLC4TKisKfMEydiCg3LpQ02OvJNElwj+CVqOPH1fB8cuoNobwIgR9HvQLtaaW43rndmTuiv
+aYHhgC7O1FYonsuwIR1AO/qC/ruNYUt4JJEXm8Wi/Srp82gvob5yvcDrE+W/lXVZJb085vjd2bw
LF7BTSIPeK0RNCPBHR4KTYaVm6Ggq4sYXmp6B74z5rzusumU/dWWlj/CVNzhOfQGUQPB8hXWDjW/
Vx70hycuc42vuUuMnLudBk4vhjb/e11T8WxR/LsA57e0+BMJlFX2NUdEj6J58Isa1wNr0sdHJkrx
ToRFY9MEaYGnnVit0TGkW4iAHX+eLtrI36JifKQ56CYt0kV8UdK3QjIK6ysTK0tpf2h+DXiq0i9c
VuRYFOoX9QpPYMygoGXEXPbJL2jNGJ4uiGfKXt+wNUGGvmlH5Lh3G774dM2Du0aRYHpNp8AqzwtT
fsYSAEK3Q7JDBIGysMtEP7nfVh/u4AHBWulNoMNlUzxQj06OvUYKOMIKSeI6y4JQysUeKllC0Isn
VMBXMVMjkyzM+uu2+cb/vjnJ9HK1wHiLespIJLePAaVhLloDyU8rm/Khz+Nln5aaFy3DaJTUrTpv
a3F923VroD6ZGar6FDSdxyjC8WWUYcz31eS7qzH/Qtlt30RYkaer9DfVMfHfnNcv5C6HFBwAZHYp
LF4RPzH5IVt8oAQ8AiOxypGOhwO+vZkzOqoUzlkC0WExdDcX9U74yFxqnPZxIPE2z9ByJc6YwxHX
SwRAvX9YfBRfQ6pQs5WAfMbKp6XCl/iC+UCnzRPSsckJWEiFBZfH0kd7SsKdI85SlJ7N7Mq6dhqo
5ZYcg1mNZM3urMNTmYqkjH4F6ypjD0CdOlhg/DeiZqWytI5qBN9zP/ohMzp4GqHmVEhC45UN9OVa
7sAdr9rk/FQpkp3gJiFmsimNadiyg4fWVItmXj7WNkMVAdrni/8taKDvCY3dSW75rM8QVBEVYsTf
Tj7fvDG8RW5vjY+BVsOPo+L1rQWKmE5QBRMVapXbLxfJV2d/1NjG94JddxfqzW3HzTt7ahUGYqtW
Sd0kVqaY89DrIz1376ZwTAD95zZiF1TdHJ8p5Z093TgAes/+JgpclF+NSTowFQazdFCAu6QAq7iP
wr0QLJ33WRgJr6+1iZ5vDhAWqn9f1bglyGDXavRVlqOxJUVEYSmPjtIELpJnW8KS6ji6qZPiASfw
W/6dBL2F/luLaWGpVWbNzPI89lMSF0VM4zFXKno/5vi+vclOkiBc1RcVDuA1WYSIXAjTvUjFtAn8
EM9HqOVlKJ3vKaYcHS4rtm4boHOvJuciQenp6EcbcWlmyNLe3Za9eYbtXfX5ortt3Xjxx5lZWoIC
eqt2AKCh4oh1a9MqGEhEzfNTYxzsJmkEoiPh7eTPukUXkDFRVod/7xCmHnuSTweRMhGs1PyN9kXW
VRL2l9hUwKXC4n3J37vdpDHKpdUsrKHagNqhP6dugcaNnG+RGD/3DWn22EjB8O2/i/FePYy87tMJ
QbLMg4RofV5gcfZtvJ7OOrCZGHgyQv/erDHy16eT5XYOLIOhSIT5KMR6SHkr565CywuthjHN+GQ2
oGWlDCxcKIWUqp8+egWsJPKQU0VJHC8QeDdNCt5yu7GffX0JwBrQ0Uox+XnTWSqaLqF8NqRfNz02
a+QUCCXzEx0HroIKoKItGp7jc5pqQuUEC7NOBmG7LioRL9nHb3yO37SbAj2sPLMsiCTCwMsTB+f2
RYis35dd3IKa+ec7jX0ccPPa4dN0r1ntkKxkS+14yvbF1E75xh3PycrHZjIkRL6bUleIDBrtqhJU
u2zEAAM0Ssl+hyJ5i2U+L53cTyKpVqdQGySmKfrAXNLTOwxLenZYeY64Zs81Dfft+3rxKwBBX6XT
z3yNz/AX22+PZh9MaIq83fSlfVkKTC1BUVDD1tUpLroLjbA4EqJt4p/sXEVlg3y8nbM4rUwoqIIS
n6tWl7IfOwDIM1dZWkndGZXd1vploLa+Wms3K2EW0t1EruYIGSnswQxHdKj+ax5wBGPMVq7UUvmH
phqmmgncbnD5f/LQCPksAX/T06xxnsSc+wumgkd0Rks1Zzug9E/O4Z5NA7pb29lwBvoDN9Dk7jTW
NnH7Z4f/zNg51BOYszoZHinzJEVM73Hv/4kA+YaCEAwHgQ0l48AU94FjQiBtf2jAm9zafq+6jZ3R
R3ETiOJ5xWh9hCzV6d7kOVyGUFTVjpI0R952a9Ye6bZaIVxVb8FsInF2lnfvafl03VID589hlQHV
TDgozXdIpKUnKHovNhyqFlcAIe7HB6ouiS9iVp3qfqRORGLjQy3HxMZL/Q4fyE5e43fGGR/6h87P
ZHGE/57C7oGtnCOSjZql0UXDUwDIlqUBNxNJ3UApzXQtiZND8B6CXyNtK8gDbPwof8xAeE7/nC3W
k9lg5Jt1ur06bWixSTmQjG7Wi+Ke0Fa7Fb9T/xPwgQ8g0PmLavCDF5wEhG4TGLYVu8sXKejlpSpc
y1Rceacb2N4A9NOePJwPt1fMQXv0ISQSX6rOu+ig+wWvV+ozjineVQM1lpWYlGemnoey7wCkYNd3
RYjPP+gWQIy0tODE3+y/BkBnkZENRYodDh21HT+9qrNChVBsptV9sP8A9ECmmoNKD3NzvPpd1LjO
tsl3e1+medzXTUATX0fwFb84+SqBJyLb99ycQ+jzfnDKFQElv/HdQoEqpU75HINc23nRvUQMeR+u
coyUzpXHnEE7e2bKakisnz7u9ks5ZXGFNz7TkiunkIEnGXDtDrb0zLb3wq6eapUyJXfRzkQsFEQD
YjnG57XKqgzsf5UBs1JyD/OVPG79Zs9XDvj4vYQRwrNmkMu4YsrJAM6HbmUbAKoEUt+/PLtDKUbM
tbIVUitlcJoVcDtivoH/0zeoHMTKriY3f5liddsZAV9l/gyfjE4+FYtwcjvEQmBlvMb1RLAtdese
XdoOjN+CeC4ZgwtSAaRkAuAA0Ylmii9DN9AjiI8vN+RYYaHge8SfNz6d9xhaRP8FnU0asOWyGFph
mD3fGO0pjguyKSCh1hEEHEMX/Zb7fOTrED3ShFPUaKw8Idt7CwyHa6xBQIXK5b/YFomuUmWd30hG
Q/vCi4+dOtE607y37k0PzGKJ09oRwK0RXXSXvO7Z1t5t2PP5mmTVbpAj5aA+2Kc8lo+YemObHZ5v
FN//+YUa1NSSb3HsEgD8nUuC/dfz53kupd9dPShinvZNug45AIivtcuTqbFcGISswz6k1ix7D/+g
DWvsICq3pr6T5h3sD/3k6bD+KXznjTWf+0NcrvJ3EcDpG+FJ59YeAfOf/5/j7SGlGVpSGmU7Y/9n
jxH11r0KZCpy+U6pCSvKkc4gT6X6nsHu/vpktt4uB5TM5XhT3dPLIU535uJcLUhP6HJBl2n9gvyY
pbaydUPlC2/89Wc1EphIHP7PE4xtRN/P5mUdnaZ5VR1QvabPRVMhhcmYZS1oPOc9Bnv7/PCV13mI
4tEWsfFBbVnFTdQa9ktG8SPR+WYxJO4PaYWuGlcgJ621KkII/9lRPeThioy7aSp/htWm0sY5AK4R
M1qC9WF+LcdbM3UrwonbN2aJG4UFedWqh4/3A1VUF0HGff/Dhxgra4aVERpHLk2gpLh8o7ivt1Uk
JaRL39UaWFgxBgXW6pJQjuRvM/RIP3zHeF4Qpx9qm/IAlAAxt1d4rf4RCpdSMVR4+BZ0O3Sp6v9p
89rJsz/lQLhLjtSBBjq/MS/hIHqWSwOws2yq1FotPiUHHD23gOrDvbyoUBTQorNnhGBubHMgeGe9
+7GDbcMzfnd4hnQ4S7sKeHFct1TlsobNnCH2DjPtMTpV4IESZdGJ4GAeZ1GfTDBHWRLpROyVn/Lv
PYeLTk31nqPr2fldByPBoctV6n6sP7tKNCrjz6UtQlkwm7lljWMrXcQj0NIEJVtERQ86d6YnZANR
G+75i/awbzVtGTjnAV2vLqAVVIglZFgrAfLydsclIILyGquYdWfeptQbmUD9JqLMjkSKcf0TFfR3
XhuL8lDYKlIl5xhnA2Ndf/tyY8c6PLJed8JahRwhymGX33ju6pFDamjVceJsfTwdIBz2XhPqRWJA
ZSORCixqmFEBLRT4rWkYM0eEigYgLEYUk2SO7FDTmlTY4ayGMPvRxWHee5XCpdwPQpOtms9036Pz
+UXsOEG1HbdvQw6w6GUA/pxwwOcmnbC5mMrqovpt+233XczL1dunwL4SWlVSl4rrGxQdpq8rpInv
xqaQ+VsxtPDatSAqc0F0VKtriRgLwrcE0PCkW+0PH1UAaRjnEPQgrzxp9ygFZAn59H+xRcR5Asp8
TJ7oo9PWvfYRvJsMRSAu7qThl/bOIYC/8mMzXblqd6Bm3nTHBnnJloj+QYyQOplfrAp+6YHLh4Me
A0HcyPwcX/neNOnwHh0N+mluHHn+X7cLas+eK/Amkm5sple+QAoRa1Fef9pF0SyQnLgROVQZ0fhr
EJn8S55pTubNeN/mNJ6pFrJuAciAyhrGPeSgldSCk3JVjx2+MiCeRr+wwJzn/FO2giegXBJtIEVK
7aonb53LTHiAEMqs8AdZuoJ2LJk97UdiS1zoQaZtR2CAYLOuQdoIkXfK0HTPoUK1WKumpVvwLYkU
rve3Mb237rwPTwjAEloMeIM5a3nky4kkoLcHG06NL34CIFfkV7T3CN8EwoN9gYwxhPQWKqHiy+mr
47VCfJeUAu1PGZwR5rvfa22vYJqMKIdSFWMym4dUR1ytdbzZpthn1Y4Uq56LnvKcFi58K0qFuT+W
bEbh5W6yk9s0uL0T8+aEKQRQZEeEpppV6FzjtA2RusVPBYL84KjNRdMzTWRLHctsdGufrAsVThAr
we5CbHaNCUPpvDz81HK53yg50mWW0pdOuP9kx3vZvY92iOflyqyGB3WqF+QCK6qsu1M/X/hBJ8fp
RXaYtVHtPdII15mGqmCUZ/EJIMRRIBc7ncvC2Xx/A7d5WkSlK1bWwinZoRU7i1/i0jcl8GRqP4uF
xRo5sGmZAclM2p6h9nag8Y631/AcQ6I7KXS8zllmWB+sLsrca98IiylF2TngJIOdplysNGYa5R04
ThR4Fu9AFtQ2xpsZLufL+ixdr5mNswsejWg0SbGuS6QI3A8QBuiDTxetzCrSx7k2z0Fyu+6L5prJ
TCl+3FfVjKm7Fe+qnchv8udoLmnVeBpXKfxAG8CE6TbPaUPX53vPbC7pm4VT4F5CMXjb9zT3h3E5
spKDLxgUch64GUZtzFORxwjXy/ZtHv7QpLLXWm6Bx/uTXoqOdJUQ4MrZD8v8sJV8YSjPmOHw53AN
hd2nJDYfpf/ibdW4GbQ4LtIvNDJ1KtVCIFP4tsa2pKYr9S1MSy793vT+GaPRStkVQiOXMI9ZjUbu
u4qZNi7wUOeLepc6NKMDy6XLg9SEFv7ANV5SBhVeg6fArn/h6BzYtLCEhBr6kqo8uXT+aEv/8QTa
9SEXMnSUnqxex/kd0gdD6jQPBaZ4CT7/5SgB2/Tfu67O3iOvllfrzlVvKKFeXdDLoa9Clq7ZvDQp
xqWUxN7XvH8wsKYZQkQcGr9EERYUQP1HmbzUc1Q+v7Bm8eSSp70gwksuZjW6HCNBYZ3QvDER8kkE
flENtjUtBA/Y1SaplqrYvvhIhAf2CEK9pZSIsCYOKikb2Hv2L8ssE83lptXSacS194a3U4xfZ0C/
xk/em9kmMYLyjVq2/RkilrCYkwYZgMgEGtA+313e/hQxiy3mmORkE/xnqpHJZ/MYvEigw1tbCBDe
Amokx+iGujPVCY7Ih2icN4PwfXb/CnuaLu6+mQ3knNryT8M+rbm5bx5qJNR97J9Vb+kOeGF2f5mg
iaVZeN9yjUOp7B8Nd25htvmLv7giqHtoF3CKUPnHoiAJYWeU7zjfeGn49SOUpxvDbpG1+ab9DBC1
9JY6HMFOn0Q3+VBDqLX2eWPsYMR12x8VAZbx5NLNsX1LcrWNWjnX4tlAYCGOHdR/ptz9G9oal6NQ
vW5FH0s9A3OIHL7hqzsETTOLEMQX8bb7NifWD+XQe3/YDEj2XHLJgYJp+zT3kwqsMkOG45SoiWUl
/iqsXeelApj9Rap4fMMNgUKjYugN7zp1vkAwQp2TuA6aL8k/O60tNH18/QxDuYCjmgwxf+hZnhxz
Sqm9Tlq6WNInqolqlEQ7cK9fQ/Z2Nwq6MP6EZN6S9ZXgkeoXTMNapan/fAj3qmO3+XUjckUgFqF3
VSssec40WLTWhBvpQ5ONz2/ICp13k51E5MZfmP7pmo/ES3ZKha61+pL3gavm9cSGIwNQiFuj4Pjj
MY72uOhPghDZ0+/h1Fsi3K9qgcXr8Ju6uRYvULRpeU+x+uJKJnEO7OJigrYi8VCGbY4ZC47VEOh1
7t7ggTyPfFD41zw5TzstC4CSlV88RRNvrZK1PyzcIa/IsPpntVwR5m1gDJOhznl6zhSZe6Cv8tzx
BYN3FpYL+baN281HIjeUatuwWqPCl+d+pHdJ78NiNRjWkU0Q+xtE1MHrNm499SaUqeRlB3/71NgD
D9EwACTfgKHOCFyyLBx/JWLQvCXyljxW1DwnVGHb0NqkkTrX+OoK1oh9z5B8XnAhYRYhOa00W0q9
TQzTwfeC4C6Ko97zlGm5AtzERL8x0Zefv6KSytMC4GT0nZtpg4OC+3B7MoHA7MjCruQ+fdogryKd
AB0nv+XPBCXQjt4YPYwsgugBFYvwFElXxwtJ4csSsda3q2ML3ZCrwOTLAhJI4ccuqBfEfOOjp/No
RVT0H2BO203NM/uziwPNlVOsFVzz+ZS+/LtgeJUgzu6fQBiOmrwo6AyP7ce/jL7P2K4irgsQBmKd
hTflsCNMaIWGVsfV1XElbFGmsfaOmJTeGZ3I9330KE3XJHRus0WdN2ofql9PBSS2uK6WT47dxdAh
S9h7KGGu3Z994djUHdPeLMl+FIjvc+i1VOnaPQBLpIVs00w3A/zyQFJXQZrJZWARmUUiGV1yT3GU
+89KWt2RbLCxZD2Pw2Pkfcsbw4j7GV7nvvozulmH/DsAfkaG9SYBiTsnnG0wxsqJPulsFUKANy9x
9DOjfiQzyeuh3sikpHdxp+TR9MMfD0JBbRXfctbGUdOskeuLPzUXkYlnm0AQ61+mbTNBxQ83r3vY
VkwzSpc5aUP3yv4wkTSGDHUGUhybU3rerGmebEw3xV5VxPcHS+xF0dXC1ajn4h4fs1WtIxPDByqE
6LcKE1lDDQsX9Eiim7LJbw194xJPNcU7kqTRxMLcSnss/MMfxkK3DBerZp6N0cufBblx/GLcppbB
oKlKvJDGtXyFzXdSGDOVrzDM3oI8ijS1PriTxhcB7F0YOvA1TUCCjMnwHQyg3DqKzrVin09Gnwjq
8T6dZT++qWca80EUheiPCvp3McqtlIpXeVmzUPROwP0uaEFIwyalK7Hhe0yHP2/1nz7xW7JOiAMy
+ON3gg7BQfW6XyfotGg9aygTHIRMijnYwc8Ng+ckNjul7fB9PRPbfVUVKTSdWIsrlLX/Z8/EMGmJ
XHRN8i/Iw+Dxm95uzadP+z+u3aLoeCOEQtEtTBVfqMOz9Yrx309nTPpEEuTp3AbkQznfaJDsGSPu
jqN0G5tzC0WN2JE4aFL6GGKYIOAi25drWAJlj9cKeMZfPRqwotF4pRCE0VaAZBMml8YPgQ0ynq5R
KHA6S8kFCLCKNWOsjnKNDiolF43l1tQZD7bfAHAwLKghZ92zwFpAREAgE8HvW3B3VWbxNrsUAuph
2JOBT4PZEPbAK0r0RhtK8GO3qEOCIl/rwRTLnfI3DBJbeoGhHsoN6qo+Uui0m9eohXcbIKYa9MaC
8kG2JGnIBSM1in58duaxcEDTkjflGuh1zZr6Ywl6nRXB6ctT+h7wBJl8qUYqlL+RD1wBhlsjhVW4
SNZeQwhMm/WveU1fWKxP43o1gEFYBgpjITKh03JqCXnz7HTgRrYIP0GmLYH1P91MFT2548FdjEt9
DnR6nOalcpQ+nysQLNcBKE4r/SgFOgI0ebMFOzl6rvQdbYeoCIKblWB7A3GS6QNlrOz9OEDZGe5u
cX2RN3zc3U7xsdmGcwFh6firBpXA6DDF0TEOLAVCLAaFtvyNceD/EMJLCuqWWQQq4wJGH4A3Lwrf
ovM7Bd5L7YRbtUiGcKoa1Tvi4GWNfef9AkQYYCC0N0ku6x+unfUdR/6k9Mn5FG9OxPImXqYfTj0/
FAmCyLEC91AKveH8o/3K32oklYuqWlyb3F2cUwWqLTnIO0epLrrOlmwF/uyuZLEyx5mGpntbfzgX
nBMZnFiMWqpNa6kZVr94eoFiwDF0vajvtcuRdGYEKdCdyc3Bj6Zo5quIBUWcU2RfMb/+II5bN0/g
ToUzbgQKl5Xz6AJLkTDaEUW2/HjkierzTo1v7BXoM3MfpxmzedPqze3ItcqjEtO5yEg0ZSc3z8W1
3QLoF+NQ4pYGr2w9osimZCe3vIh8UcTFzWOdt61CoqUX7JdSJjolOAb3TZr69vVhMXP61USXQEB+
ZD0eIO46nLBgJ6AjNf9swIka2w83fvMMu7AWgJZY8rhS8IKhu9LHUbvUPmwDXw/yNcGNICJvkgp4
BH6j0J4hmcvLHnyqoTNVba5UFSQL1G/SDHJURnHUKA3n++ADdlKaMw/yxk9rBvZINPPFed1rhLja
EjYJfEZsIJq4v2m5bE5fOD7P1mNJDoxEWn0scVenvDrj4YMM5a7WWtgYfrs3iKO50Gh+80SKsJE+
LQzbJR7YlqnDlsBqOG/qv4QsRPSuumsCqIzMAKSwTh08C82WWejrS77IeJu8b6Ds/kF+KRs0HQmB
4+g1Pc37Jjgy986VlQ3UvNCVRtjlpeqEfVY9WYkHIVnN1SbT7kRykt3dD0VwnvENqaIxMfVwg58r
lU55973uCt2vnSGND/Wnqscbn8Y7j0Xa2OHElVO7GIF0bhVTgBdhUe4dvPcfGHUwYZSGZ9SynSeU
YqKL72IYB/bekijoaVsxsaMFxsCTl+PoWDqvXe+eFQGB8GKXpzNbrTs0cEXJZkzIwq57md/R603H
6h+g49/lFZ0h02/3I94YiFZauIiu5J/9wMN3jLYc52pGq5jMivfa0DeVqLJxNAUWei2haFSXINSU
TgIeLVohujBnQn1GFfRMLps6T2E6fIolyG9rpjlO54oL5o+lN6YxLfcJNeaq+RZUJl5n99+PGaEo
Z6TUJpdmEtdH+obVcjMGiiizWGIc1G3yNUY+TASUGJytjfrNyUBbI9F4KnofFvHvhyk4peKnNzZ5
FnYmwBgtqF39gdmwYQl9odEl1WL/cafVx3CmJ0xlMMsCIvHccS8/7HPhCnvlzsnfZVCptuLEJCDm
/urJwEiprKJdNEkplFqpykhzPVjcK7rB1eA09mjwn97gZhE3SyPSYi3pQG3OeZPEil6YlaieKufR
sWRlgzq67gAG22KZr1g6JUjHTIDQIuyTZxTKnCutYehSKUQoztBQrHcY0fyQtP/NrdTrqyXnu4iY
ZugPcoP759TpLFjYbS6DLxESdNovoeXldUe+ZLfEEMC9TP1fIAxcX/ygAgoLIKqZ+i2hLuDBIwz7
YgPD+e/+GeLSk+XH/H1lnGVMubuEo5XmDbvJPjpr4euPiD3LgPpb+BXr+ryHyayDB5b9Ku3TQlNY
YABZ8VMLuWV1AQsoBjTRL0tdw6J7Pa5LGBDDQZ0xNCTtp7oj7uXphgc0auCnp6yntHZ5omigoqSg
NqMhxN5lZKs4gS7GRsELtKLodgb8mUvouHPQPSvOMLnuh16GAj8E0fKwqrR7Oyvx9krCB10h5g4H
2zgmbyj4NmfpJ9LEM5zgErbJqOH+d3R837hLR9fxEQb8WjHMtOpHjkjHgN/3iO6lPbnzbd+nM83i
7nfOwI8L/UM84IBapodDZADZf/mV7iCReqtfuD+/LpLe0d5JoeWBynazDeEOnwE2nIQYxMjd4DeZ
TZygl+IjSrC+dLlaNxEQrXLGfVmhY9/qdjerK4lqxySi8X1+GzaLyFjMhipPVPiLXqAYXVdN+XWp
qBopt8+VZVQszuRNG+vPl7ev01XtT3JYh5wgxksljE00lW+MMe+Vyiwx+yrgPF0iVQ9RUKZ/P8gZ
tZcs3vFR7ypQZSCpQSLIK4q/AWpWVc2gUSvk/M/ulDwt6TCvSjIGzmz4Bx3LPop0JOR+ihPalW1n
gkcamlYmQSdlw8tL97WD8CiznuA47+qI3TMQPtD6fhlPVg60jS5sxqS/ViCRqxmZuef3KIhCZRyW
3qhFHKB+MYJ8LWhvatysgzpXeM7ctMXddCUAZ06VpcgfTrpfkoF3e93PitRAU+HRJ7tsqGe2h/7+
ljDKgLfYlwyHNtgBhWDyv98Y/ctQTsCx/sQqbbY49yo9YbvvyDfOaWCDfbK/hEiD+h1Sa7J+xrDk
CDm338n3+Gx6OWTx6JuJHTvmjgeX3rXMHbFQRwy3lvJDixvH9U4IaC8GdDkUjAazSyLbC6/O6Me+
bbLgFFGcT/tVMlpzpXbZhQ7v2W+VK43E9N3MluTBqn5sI35L/DDCm91HE7B7gZhPpGbjv00j+xg4
vLUX0KVN9LvxtZfkDKX8C3D0RauR+gDoMmt93ww9dt8Txzqwto1aujcV72s1zEveN1nHZGbEJlnI
a57FRt77xY5VSSMOgp2IOd0+Zx7Div5w1FkaHlcBlDhamuXJWdaU2F3PyQHJGTVqvp+m0P5uehKu
Z1P0KLYXjAPWueCTNCFkpUii5klTSYPHek2D+PEjbtswyiAKgrqvwPFMEsq2S5EUnBZeKWXHV96J
Z72iSYfPrGjMyGtg+nCEesOuEre5yqvaM+6IuRuRho5Azc5okK2umAuQVUBYe9X/0Icrf75TaLoR
3cN6pCrBSJVc8pw5EDEEnAlsqx0P2kZjsEziSLj4Ib+PGsk/kmf/DDjrVCanggLoQXuVQRscYlIn
raru1MRr1TWTB9qTbWF2NR/6Pbj/PlPPawPdQNZ7adPRgx6+5Qk1CS5rM9SYWBeMecIdNEKPWS43
evBTsyNINjwa8ZMj6qkHF9PJHUIZchcUPkrP3dr4H4iUxhQyYSjoW7BHfIKIHJWnVSo0u9liGsbE
0HeU4K9agEVjvIWM3802qw5XegbP07uFdabt77aKEneNa8k3o1ghgsaqJQpBuqBlAG/LCj5eXq36
S3dcHtm1fsB7MVrDSDfrOUFu9Xes4w8D4VtykzEplc06n5n7D7qINu7bOTlhKrnJk3KM8V97YvOs
JstcOglQJeDowbyFGM80PrGj6uCxmqHKvlVir9QryFVekmkZ8LITp+zbah4KSos6WgHS1kLNQqQN
NySEMlVPunO+2nxNAbRafou23ksmBoxiQlJGbWBFlSlaRrm2s7bCptSDOeWnX/B/3nc3ixR5R8/F
ZoDEWw/2hFf8LYMZo0g8DKW4rKW53GWGkHPfb0NLptBzdlVY7xprhO4fcrqQg/DLwA/Vy6MRGY9t
o3xVHH1FUbBRAD6QIp3L8VeQFGu47HNpy3MCVzThgyl7GlwdrM7JgWRxXjHSgOgWfdBt6HFvF/jd
ko8CN/MSe4wwzCrquTeRm2gN+s2mYI/+WBIYQy6Y5BfSNBpgBkKW+pNSwamIEMKVvK0LTqc+SmBQ
8/tnOnQYguI3WA76526lAq5Cd0eNMcn+JTTa49tzp+35RQpMnr88YHnWegUGGnKrW2j93u8eVEQc
J18hpnYxlwZEuBm4M9Z7/s+pwmP1oc2rCaVDadhihlx1EoYHL+rg6E9zjAPJ+xxOsiWQVRADDKYu
FZvdlbl59ZxauVK3eh4BdbxWrJwXNtNJXyQvx6xlP4xMpvJ+DYdjt9BDQ21hDAzLfJHnmQTcJbyS
jOtyigY1HkTkcqQEdTTtXaWQdhDZo1gQ6pbOnNrvFQqLlMMgnRJhNxdr1j4vTsLlpISwdE9te2bW
THaj0dJnIqJnnWhZfbj2tVp4jJYbtZXDI7hm7iIifguDmegJIsbQF0HX65ti2uG7XCaYVPYA+CoD
LxuWqBdfqNYemrzSBUfjKYHnDh9twr7IhDAJubN4OVtb4o8SJXfWteU1nzrEOKA7QIx6FxXJpMJf
952tFOkP/MWn8h8dMfNAVsJUt0/Fn2u5tzJiRCsfX51u87WINOySppkg7dnntlP3VJhv/szoxHHG
LAzYU2XEkW8d52UD7u+yU4xnKZpcEJhatRv49hLAvfPOdNkc6LhIw574labNdUB3mnnOIKs9X5zI
5Ty/Aync9PWnpaQGxVOyImWZ9Wpk9A0uFjNN6g4CiBZZ7u7OrFU2eHySBvgEIC7m6/cVhDx3t86y
Bqw4FT+cOxx++OAolBgeT8Xq4plSQoXu/mJ1lI/Hb+zOkwDd9RGAF4aXAUWsrj1779H5yGH9uuD9
eEutyHQ1YxzTgRv6onPQjV6ghlitMs8vBOUbQOkAWXH6tZytAqaSKpqvs3Rs/KVjZ4XLlgLPa2Gg
BWhgDGmjxpPeANdLYNd26JH9OObAm8XdsU8+jYat3J/wdJGO5M09ZWHCkMJ25IyEzxb9LHaAJiEK
Sj1rDIHNPdfPcgPzmYK7jv38IVBTm8xOUnZMeXQ9uSEDUKfVY8dS+ODl5Dj1iKFaMDxSh6fdBWfN
SyIHC00llelv7EnQHsPhg6sxreB+sdE9mFQCyVu8QSLd9MKSZ4ANE++esl2FY2dRjnHge3e9cYUk
ZhOMML9GQo98XUApZlE6JnBDkXaXhvJ9vR7eJCAMtzYDV7601K4xqohwDi7JWKs7F487QPTYtWvq
tAMRo7xlwm9OsF3WsNy5y2pbbe9zl5TqlVnN1TZE56//Z5A4V0kACQ117Ncwg0SkWv+uB7RV/efX
eBLiXXIWD22Qo/PrQHqqJ8Q+4CIdnAazlPXyHb2KWAiIk2J9XKdb0Sj3GihlueAH9xg3le2CXhfF
B59I6Sseml4zwOOnqOnelLPwqzx3mg/lC77hOXHudUrZ+YXTLaVCi5p0GEqGnhfJPQF3VRFrxKwg
wDsA1j/h09s0Osb+NKlbebVpeJJt18UF/9jOEeD3SjBPevwGzItrAABOEJ+U/vBk0HCIWJGXmSFl
JPCucleF2RcozKnb+1DUJ4TslDonPCyu9gP0JRCSaXZO/PMoDPxA2oG+z9gu4ag6u+XfLbbkEwmO
58yHcwZjPz+EiBAj44rHSM9uQJmrGchqu6M698Wm/XZCTURDbp0Qlo9lLzocyfkVofWyQqFV4kaH
mTxh5NjTx6Dw0fEQgo4yPWIhEwu5XWHXiSzpYSsas4A7j34o7Io5axTt5CjTBdxRnB0QbzgLYDbQ
Xc+ELupi1WwvfC5yM6aG/El71Qkw/Se4OUWNn6yw0ehXZ6OJwbp6Ha2DZJBvNG9GXvK6WlpszN2v
Y8dntf8sSIojjMc32wOZKLljBKsqW65MVCQrTIcAb+Mq0QTjUuVZmJx0+ZfZlwXktPmmCy3zr90I
JFN0tPZjLdZSNHlmmhmWAAcTuBOPgR68mIOor7A6SBnQOJxKr+mfSEHgD2y2ckXhJCnBP59opLk/
fMvvqy86Rcj3tnBZUky5q4c2sqgxreHdwnVgI8hmi+AtE7lNrR4iRu1JJ4hGIXZSIGTISeB0L6Tt
JTJMgQkrN1NJgmHcUCLE17zKlUHHpysWUPGIskSMOssUuq9kqfTaxj3d3sLK/jZfPwfNLkgHg6Xp
gkbxepLXMg6RXkue+W2jzIF8c6Sm2oUE+S14e3WIZ/ne8VjiasCgQTuRTX79wR7FcjNZz7KWr+lo
f/WNNEuZQcI4b5iQOcfWtfKANtc0RvUvdAGXl8a5PMyhmLLWpXPe6JZsd/H+62239NKyzQy+iBCT
ZU2W1lN78VGebfPU9RASxepd3OcmgtgIHNG7oiZFb+bq0nTkTvZMb0h71+4N7eHtLswOtpnKiCKb
TaHJ4ESK61srKgj4u6/+mnupyMUf6IcByRwFQugEuqi1rmAET+muAbRw11RuAQv4sKEbXoI8O1S2
TTm/G7FTGUOHcA5iIIPwrKWFXaqpvlvDekf1TtAsiWsM9II/pJPEIp6VCNbSv8lRBmRGMshjXejE
ZRY0hc1bh+a9xT8vcQq9chnCCQjqmhXxAxefEVv8c5aNjGmVLxgvvOzPGBhZhdQdBc+d/ZJLajdk
L3pZkPr5di5iB0NoHoT0holajffqD6w0U/3hMzqVmiJgaqhs4WF2n3dZu5/wajx/8l0teii8jPfo
xeo4gkA5eVCQ9rfTiDUsHPRMOosgvvQjC6yAH9SjxTzvJnzHLoBvXbpPkUkpBFpztqKtJIGDSwQZ
2g3pX3X6D6ypKd3tFEJOXBklXKyuP4td1P3aOVWT34JEgRrybLLD5PWINsCf5PqCnp1q7rJ39PhT
tDXTkLNGT6HFmHczz4ei2XdT+R4syoxvA+qyHnbQKyvrwIr7y35zkeOt5gwnhfMWFknTjjXtBTkF
IhurJNBAfw6QzwyVmhpbL5y7ND/+iPJLd+SoD4snemscqZNeAJxqkWnLJ9Nw7yK2vB33twpbZBiB
n5IjTOYmPAvrUVmSfd+RIoCt/cKH4V6z2eupM+c68xMfTGaidFhCodBjf6guLJI63m13/vnrRSTO
ImeTsEMjlfqT4eocC40B8Hr66nJ/PbaWr+HQjy67ePbp921fyqZ4pnq1vN4KonkAZPa9n7B+O7KG
OjTrLkRDH0IgVmA8plJfC8d7ehbUd64lt5yxliDn+3AhOYZfzVxmUJJkBdVQ//G6P0afYotMqx1g
YTyY4PiZ2M0f73D0f/AiMR0FtpnVcbuKtzmqYz/ilZce/ZmixTO7Y/Em/AQvvfvf1T/QYK8I9hcS
SnMon8kuBP+gFGw62sRNy1pjHjuCSiHNfdHXq7ug2S3/jVQ3b2VKpcmzuK3+Fwqlc6siHmv+oEII
6k8f5UpF+j6CzE0MwUrxoU/JvNnC+0WB3R9srY/cmlNQOvwI50Ae0FOHJmf4w1r27ffb2nOLaL3u
l3W1stv6lnpJlgVhl05UcbneaMV32sak316CZbo6rirejj/Gzjp7UhSbmG0MLqWCns3xVRr/es3C
NC99QcFnr9hMHS1bNqtvY+dVUSppw4M6jjpSmW03He5MbUWpNNtGzKYqEsGShy1IEmrpph6UnAv8
KQNmhEKzNCqvQ0SEfcK0GN3JNt+/Mp+kQE4YlFX9FDqtfGZGAYcYPgQnV1YnWtcELVSVg6Ov233w
rk3GXjaNViCbdoNIQB/i2nNeKgRWEROCz38X9lsBaWNtZPTdoFuo5LWGIkKrgIa7IrRWGGtAmjPn
UcfvmLMic3enxsNOm6kZHLotUJtMjoZi2RPUVSz9lDywmNNIJlCNqG2J+z6pdBm2+TA6arv6pLy2
LYlYyvMMstBaIIhT3AGToi3ff3qO1GVJxZqD99ZuNLssm/Av1qy7quoS6hW6SPTtn+ot4qUdEkN8
VgtubkxLCQ+PXlcmLIEUnMiYBXCRfyiUX8LcbSH6bkToNgHx3aeMxfo/0Tp3/g+kiRlq8iYBE1eS
hhyJ26vYyqfzYM23wEkZZN1KFubSXaQ2XCEK4bHp2gEnLO+xkuSR8lW3qrFADy7LjhLKJyosved2
eVerkfx5aJO1pi5KTNtzoshCVJYVqX5Rv1l1BX4EYpcFRtrPs9nT3yoJU4CrTtTNfF8p+KpUrTl+
NeOhTei2gsQ4iXjlJGcQ2UmtQNdUNGzE6wd24gsz4Xzvr1AYSUOGurUq0uqitsSrVutFV3LY3IjR
r79bm3dVMauOh1/Z/loMAXuG4R3KvNMpOqKV8Gb5dxcV4iKffRXSXrAjznQA27M3N/HBTv2EImKw
rE3HSJ/IXLoUXWp7gD5t6IFilhLeSpzfRB3F2WvVCALBF25SQBRYqlpflfnAvewE4Tz6GQgb/ARS
mdv5jli7MsumcqyLIbWztPUf5r5QLzESdlS2/Hka3FopmuKbGYnnMYk6P7JLkmIWDIm48KScqfxo
iNO7voM+K1/kRiY4oyumKNrcPGo510STPKdyFwe0sSlpUkQHLUVtCoiPOys2FyykWjWUhEUnjpOP
RBpPF1eZv2jE+8+D3FJl13Pz9/XX8r3b+btQ3URgSrROfO3LLwzfT+SpQvkezD8BYbrQjnqNmCB+
A2RT4VVgNhPCJT11Bgmq12j5vcDKQ2S2MwY6yvLZMlQSx2CzSixLg711ELEVg7virpAypZi5brha
esL3ScSUBMgDABDznbD5aTAQuxHRJlaq5dj21usyj6wAsv3nFslpaZlIvu3rJg3PvQ33OLehB+Jc
eJFWCqXa92PRFTxQLjtgYsdcNTsJATBSIhYatizS2jSGmhCJcCb9rAemddiJ9zSrE0u8l91xQVNl
+huPx1FZHaA8QywAgT92SwzcecXxl44mOcMomH1nQsupJlBYp+zIZdtJN6Zzrj+JnsFsed88bXJ2
fJ4w2zcFwlLzhd85kD+cdzbw+n5dA1SxiLDaT9Wz/qt7TbUgegg7tEOXIzPZAvALrp9AYB7xnrjp
am6ac3LESaNryK2ATm0NDHO9DM8UPA7jpdyEyx05WUCswuzIv4bUqZQ3oMncb52a/wk3pxwMdHqY
7h2Eqxa+LeBD9yveEpp4dwGwHTMMo4EYgqLnyYqlNPm/fYclLslckpz636nx2v/fCO41jYoP13kk
FseEGKKhgSizqZCaTiMaYuSgZWtOcz+0OlGEyJ/lqEDTUTLfcMn4IfoBsMHbAQ7l3wrxPqtd0aWX
v6BPnSWcx5qrLf5HQ+dPvEWONY3OgrS+CFah/df40rTdEo6W/SE6F1TBZzsJJSSX6MwxJy4m6In9
NOL73O5wvBdA9EGtkxUB8m9P4onSkLEhaI3ZrqYzDY5jGE5SMBOjkf/I03brl3tv8x0fURUA5HW2
E1XbNpULUTPQf0sKE10jwcY68AhgPl8OZ5iBRZTdhD/EMtwOQwDR6H5v9tEM4MfDqa00USMUJa2i
/JszJloAtqrFV159oDnmOU2ALRCTrasBLOVXUnn6+IR3ysrtMqWgT3dqvCVIoZPeIM3f9xHfvUGr
+xqH5yth4iswbwcciiP5zNymFtzLAxAOhq417cs0n1KjRGfYciQRXZvXpg0tPt4bBE+6H+umyiKh
Ib2Zb0PHfQWYn6xExUlUFM0rDixDrNKr2vKSqtFx6RtPRgFnzcZ/xyklArPM1Dn8BpKMb13N+OuR
oWP1dK/FE88vUf43WWiSvQao3xYoe0F0SLeMBPBCd2Rrncro6KEJUn8UiZZeliCfl/3DkPw4ykmt
KS+z2QiybuY5/5qhN0PMyUEDu8mthRGxIhLZ/L4Pnsv8Ssw6KdotRRl2tTQj5kTbEOZSvslPkdit
82hcGBuTFsrJ4MhNKRf32X1tDdZkV0JQaK4Fuxx90mi0tHLcecZyvl5rZVZPQVf/TVrtRyaTPt78
JpaT47VdGa4rOkiMDKw4OZE32jD58MRusSmpfiDg73MFHNsk6cLmcJgE1PnBp5e2SZlPVdPmMbF6
Xw5wuy+vhp5LBop63Gm0yJszmkj+RJJ0j3DBXc+lSDQEORfS6GwF14XMmhAM6WXAhkpuLAL0H3vF
lFdafmzjodFCBYvGXKm9w3RGDRwJT/RGxW2g/+d2SbsrsqqFCyJiMcSR5MJd5iEmgGqkQR84sSue
Z2/Rdsnu70ofJEiw5D5yOOtRUSJSPn1FzKtuagMkNHVibivma2If58HYAqn+mnNZEtfFutjFPsAg
QQ70l+WVixaa6ymzzbPv4FWG5a/FiI2HIkOU9vp6o9jpDgyzPPirdnsPfzd/7BQ+y4nS6KuuP4N/
CRmFQZXbtJfXQG3W/ks44yzdNXKX8uOlhNC72593XKEJzYFf/I/15NL0DJFF/cuoZTa9LIr1TmhF
RkABC+n9Xt9j7n03HZ9QGHKDAtRXGqoo+G52XCHIId5L1yY2grDrhi4lz91+tEhJViMiXbolzrNa
0mZYRg5/btura5AW5a/+tdRG0/Mui7uDodwATHeG/bOuLFg0J1jJNsTyCq2Cppu3bLaYi+kJUXWk
0CCgPwmbZ3zn0ABSoYSAa3dFyNqL89yADOHge0Xq1sOamWpWjHqwuVMSITgLYKK94IbWZIL5MnBX
M4ErMelTxFJtSvtrhBQTiHWlJk1/6UHbL+p7qQV3WAfEoF41yDgnhhjcTq9N/wc3CaWms9ucuRlS
dGrihD+yZhNtj5mOkGl4G5IsADLUjYAjm1Qj8w2GbEpUm2lGNVG5qJWiEoj+w22OBv90g7iVq/0y
A5/EYUFRlGgJuWPEH1atXZ8NEfyU4xd5jk4qvDGudnu7w8jv1iP6EwxKt3LFZcMbcGne4ZoT1ukl
uaK91cfbpIAioFp60DEAqWE/JB7tsHTk5SfLY9Dw1Wx9SwoA9ygpxTGkC70xmT01MFs7ffWNGUTD
fSzj5PI7wld5BjeZnSji+qcWQ59OnLp461FI3KQq0wCSs8IKaOoh1dPFDmp6XLzd2CBVDMO8t1bA
L30vfvuIodkkqb/4XBm/GdYPU/F14QOdq+qzfdVC8NV20d3Xdi2qfGjjPipmodAuFI3U9n0ndOAD
sQaH+ZASOYi1Qo0PJdkzPLz2VRZ6r6MjJuxvF3ivGcv1uNuPMJzQuKJoutP/YpEgtHNMUJFIDWVh
4ZlKmarzU6zn0XbHrlUr/ZpBaDbspjHNOr9XFK9JPJDlNm4XlTum2s7Yy3F0ildPJ/vFKaGZr7fF
lfi2XsNL3lUY6CpcSBUXgZo2S4/SIST3nFvMvlmbuE6yDjx8KQpYizgmggkuVnA3HmAAAuZrQHg5
TRJhUT6t6Xb4p5Q0z0HgKltEqITwXbNI5HeG0FLCDs5Li1Nuxqy5SEZAJxzLVyQqGoFhfc27byKf
UxWxBRRFe1wwkfYu6qYUco22gCZaboT/kvhkiMkEeBDv3H3jUje5AMSH3Si2oXEZK/u2G+MpWuBM
3lwyLZB66W+jJO1NlO1Z9fBhah5qqjJcy0LUEHNonTqggJavlO20n7pVsLm5ETJd1D0N95DPE5GP
J92CIMzaTTLvBc5LPtGjuyvgJdyH6feB7937bU1zxnpscxsqRj6a+fpWYfoFPvjY5POHWsOrnBjT
PyEzEHqSthSnTpqzfoqNkU28NV22VPbJfteonF3xZW2ZbRQlFd9i15NKzd2DyyesdQU2LNLkexO0
MONRzipy8nBlXxcaGtoGMZmNDox8FUZB0lB1iWG+afIPyo8ojXee2Ygti/jFHvasfhc0Ba1D8o5x
q4kjxHL3krdaAhHfXK1JyEXOoqfgL6AbUMhbKKw53qCgxHA8KCQvozhyi3c1VROInq8PzaozuAUK
lqsS5qC5/9ujWzvr8n8ZpePpG55mVABmUqW+keSdCIFIhPsYBbe2dXNK6LBOcAVcdsT754Vv0DI/
6jXe6AbdeZHZTlXC8JZH4pT4HLctF5LBZObJmzxzj52O4YsFjS8WYj/0OsMXy0501XU02ek5mxGL
oJyP6cyXYaaObWLWbLF2TjqzjVYF/hUatzDBgRBcvBbOESfDcCYG65u3M1CDwC/ILOpR9T6mbIS+
8WRZmBWxyVJ2KVLGA03FncJcPNbxEv9N8Yy80eN+IH4jDHCRSnyzRDwI13iGrdiiukXmJMHX7cSE
Yg4LArs8VSXYjzZCk++1R6Y2sQPeHwjQpWuP0BfGIMhwYaCp+5W0ayMsYpnmiS9mfAj967UzHnsX
+oaAVg2LYdz/PngQG/Miv32VpbeXGyL/gYkSXnE1AftOZBppYTHD4ivu8g7MnMSVvQ4nNTO2bb6n
i09fV9zBJTnR6wMMhyJ6eP17QVAPNYmZhexuPvUMzdcixmixqqOZrXXYzLJCpF+mbOxUf4Od21Bb
sJ6SKW7BAbcejhY81yLWrhlGoFHqU4hUYxWGWRcdW9z2F1GwdXB4s0bA3yTxZAjmryxaoJUdqwiK
Qi5nThhCWCZ5C901iHZDfcUK26IjGlHKUdz39IaE0bnaJQ6hqJBDBl9quk1d4fdXc0sOuHOMpGu6
5El4ahJJExbahVSvuT43g6/v5Q2LfCbuy4Bp8yfUFIy3vTwi7cBbnTaMk/UVL1CptixJithWJUCn
WPMcEImcLKKZpTjBfdDSkyRv1A2jSaO27AqEQvbaGS2SJOhtzmf5jV57bbMMZYjzNpd47Mj3C8/k
VNUv/u0dhj7eJ7YJT+AhySdx6VV4602Ptxi8JSziwJnygURU5xLm4l2ubyn6jMc1rmazUVJc4df5
jeiZljU82D6gu3lnauYsQ4YFa3lEu5ZBUKGvyTSrFEl0jd10LHqPGiSs6hAuHmQSyW/4HxQwWJPf
1QwyRf6NedlozqdCYKXVqpDqJpyDx36haTgv0rCUrNf7WeJvbcbLJQyRlszsFg1hzfK0tBS3kGb0
v//gzyO7PUWCPuq3tI0Rn3hxAwhqPL27BfbPxQ+VNIKiUnAe7phZ3YNiz2rBOiB5OA+zmf1j2Skf
0Dmb+E79+kFhEWFuvY8eeTepG7rbhbQsRmONLg7wxQXX1FtJdn7TzVJbb/GRYaHiaQiykf+1aL2H
ESXICtiMeZ1JtGae985Q9P6jdOcJQehaSlkmtaxcaX/Wu/I7p1o1etWWf9BAIirweKlbvaWXeXRE
ceOW2z6kty7JTCHKtXT5/RT6vFgmryQCiKO9vlO6QX+gO7432mAZnjPrryAma+WbZEIxsDgyUjRy
avUqdw7l7gFC+8C9/mS3XcUR6oGPbK++lRGCqHRYu6Cy4xi3e5+DPXaEDDEOvpw3BiNt048aepSN
aR+HjXM2s4N8obMAzvQ3/xg+1ShS0rk1MQBKDlWYbGiJ03Yztzq3dgzeWJZRbjyF37pu+O3Ob7JI
lUmFnAaKjutG8anGR0knTms7VHq9nR7TGcZGDwq8hM9USladH3FATEJjznL0ZeIu5641YJi2ZTmM
G/WHFxcN/C7BnwB+UiQycbdpoW8Lz2BPzqjjqL+Gt7QjjJZC+kTQXkGFewR4pAvU3435lCto2JOh
HGFvAjjivXxqfOuWkfOcZvuK3XeOU/qjAPhB8yJMgZXTmPo3I08qPSIb+htgTJBnYS+DGqWVwe48
khffSWHMBASoGgQ2HIOLXFuGdg+ayA62lvZQN/ioZ5Yk2L/YxotErq2cXi+NlHe9JfWIqMea+/ZY
9hft8o5E0UuS4fyqFypzqlJ5iG+0T6sOpVwpjS7EVVuQJ64mAaH7Za25Y1iitVptIJrh3PR5V9uQ
kCLPZYPEUsWYkExJEgAub+ma5sZWgIfgrlMfsy+gSKQcDerOeUZ2s0UTJsUGLPyqAw3nubYdEcOs
aLavzwUxwwx0QhaQRaJmOXrp+toJe0fKdSp4icWYsvQ1uHnigIH1vbKGMyjN2TOvqOtJ41iG+mo3
WWcvB5JhLAfk80K3wFpfWR85h4DO2MOx0ZiC6CjbmtPaWYG8iDilmmA6dS5hG3+IXoLBM9CJHq25
UJEOPvTpjFqX8Ynq6JSAa3MoxWta9UBt8Aplei4ZteXUESR4Hb7xe4iQQYTPeD3WD5kcR1k8rmer
dfVt1JScFSpUOP6B/k4YFQaSbumQwAH+Gp3dbyAfjEaWm30xQih+pPdgtUOUifQSDYL9DJeEDTUH
H0u4bcpNOEG+PNzM3zoz3WGZljLgMEDslkX49iAXnQOLuETTw2fc9lFa0nvufCZ4FQzLfSX0wqcJ
69bEXl/KLHEivv6dpogzpRHaFdOpAhGbEhGnmkVD8TKENteziDS7qyQwvd1QHOHZ6OhlkE6fzkKT
kHElHKr5Zx1+V4Qexk0d4SQ3OwXqYP+lZVmVLkwHCVrfmgj0X0WZ2P/N7Rjzv7Nw/NCOwGvWCds2
7ejBbIxU4rnp0mEYoDpk+wgB5vBhV7RLsB4vzgtjc1k4cPNrFwuuEsKtFp4+fLQ9f5izmUAiuPuj
EQEs2SGLZHESynEr5BVQEeo1m51bxqpjcBcle9NcyxjX1fbDd9DEffyMC1hB9eASvsltIKmc/Wjv
iLpnxBMGpm0ldsfrPVEJUHnObbPlUsGdazYm8v3Yg0QOgBq+0xeFW3uWFYZ7yBVnDZQzcACvySX7
4+pkoaGBLZWsjL20kdRXCAr1G/ezThBW4exoDBQsDaInwcUpA0rnsZZiBtu5+CectmGRBPLA9qI0
xqxX24MmpyeqPpy8jcV0ish1V5pwJm40DFBpo7biTaXIwVv5eyyQmxJX3jGyyV6uzizJnH0g1eg7
RN+cBVbnO2/dmKpt6DoJZPHSXl6qTPa3SmK6b0YtMou+y+tGsy290lVAlZqkpgMHQ2N/1aEjcIvq
N5mGR9x1Q2xSYhGBlnIGtcepOnv/C9NwtnP6lr0yHs/+/uUmd2fvFshl90ZIo7r3PrBRb/TQJzR1
tu8OHl3xEljd9RoQJBYIG7hYgXrW1oDazGq2XisVeYXI6/jhn8IyRN8jyIl8xb2A9B6fVWcZOQo2
HTs/0H2p+jUOc4pr3X2tZWhtohmWEZfpaMh4aPIrtJmLktMfkDJnsyOBKkNdx3r0XKLBp1FRKMXE
wvPTP1tVEJ/+enhTYYBBjMYvSITnVETDcb1MHHR3RpriNISn9dJZ8CNrh3psS+Jd909FiDgRqfW4
FWqFbEEn1vQVCIfkO1FyPdsok59RROZMfjHdPIwdkMrbKmQnn6teYrnuNgefTN00nr1fU/JrP2Yc
maw4/Iz5bcVz2CnU7bf/Bx96HPrl1Knxli8nyrGcSaaEv5wqicpl9gvbbIEhbUvpdARnkUqxyegH
tOpjcoihXtP8unNsOejqX5dj1b/eykEM6P8Q7bueWBIFjjXLGy3CfLZT+SK3tnRGNwXostxAA61N
aGotJJ07TTOtcetEWUKL+UO1Tbq0o9qBcH7WPgoPBjFkTsVLa8o85odwudjdCeV7SxndsoVIZ5rI
KsumO/OD5OgoMM7fWGwdR9dLDeSEuJW0wKoDWmcnrT+tOslgnKbFZDt63SItdZyCKolK43V5I6iN
K28YGrqdn7yCUSFfoVPkI0VwYxnPH3YoPr52zc5d55SbxIwO5J3sYH31xFz5fKQMnYoJSLBorM/w
W9Tn0t6NG4+9E3DI7Fkz33LSX44knx3UQ3pgADda2mmB6KFzDx4we5luqhycB6PFvEaATqjBxPS5
Cc5fF5jILOGuXR5Hc4TGPaHUgZyr8xpkT0PHOo35Ijg0w7mjwatD8Bh7Nk8p+t41FnzLJOs393ym
zGeLQI3/58b/O7zXmDMdSBlA4aPC7SDv3b5bBRBSQ4w2xFDTQsbPSeqjbTOO4BchViteGP+rE4s8
tjQ6JimtKN1wN1NNSxtM2mmjUxjZsmB2DFPuX4tTXCjBXrPGhrcBnBZcbEYhRhMA5/YmtbSSELAS
aag1LSrEfDfk14mrDH6gTZiXxLRzoJ8Oo2IDKPUT9cKoT/RlPn8EiZh+KIjQTFhuNSe8ynmSNBkW
AcmcAEMr2ZnFIzHN1oGFdu3CQnDfuZtL3cHgj2ayJdoC21Qx7lgwXnLMa+v5cUwu50n9ORQwR9lj
fNbqks4eiVVIl227OUUQxagu9gVJKdln0O/8UMdu0dCo1h9jD7ReY0VIV1s6KVxELakaT/5bkvZL
iHo1sRjmqVNpnxWNFZ0zK/f9Rgey9fC7r9m84VPDxh2IUsvIV3M2+nbZiECUIekMjZS8+TBFW48S
Tej+HW8CbDibN3i6WZyF7Wr8SaycM3b7ACyRhsw45KvwR3pfewO4NC90ZUU1j3x9rMuHNJPKunCd
1K+J+QWA4LgWb/23spUzMN1Ijjv1aDJaB+hyC1sm4MMDqwombd3iQpqHiAjCkFHutczH41ghbYhf
HUTdgD+R/Oz0Npy4LAWZGJ0qFnT8ZcUMVoLz5K4g9FIN2Q5hZE2jwSryJm+RsIhPFm4sOTHsQ6gS
4DMdCh6J11tUWGpU3vJfv9EMJJz0pdr8c8sKbSGxNMwdAGL5bomCHltkhtRVaobmNzUVcj29elUj
tbyv9PEMW6+mnnefrp8MHyzKkBgb/+bIuoBeWEOfF68z49qG8so8MBh/AnVI21cotPz3qFSeKiCz
wK5/5cF5/VTemWuTHuOuWd12juK7DK81tb5OZ8CetZm1la6kfxGZWWCACu+JQwETzYiWFVGm6KJ9
ov/eDsweEc3AF0Z1p/E9hWgbqin+Zl70hL1n9ic7WzJdHzfumTQ4m0i2ET6CHVK2d/N3ig24Motz
oyKJsJdF4JtKyIdNFbNyXGcla+3LRBE1XWmk6rDC7YPYwjp/ojAU7AjNOsLk1Mr7LxLTg8YQwlGd
RA6XrvbeA+lYRhRB2ap9FLoWsKDKCp+k+NhXeLdBiYor1lUuFTuwzXtx1XzneoY1/nJMza7tT963
I2QArFwKrit49ZFezwy3JxFQNnB2J3ZiS5Gb1nDARttONZvUZVTIyDpcxFfACC3j2s5J1X9lwKtx
ZUMNwfqxZJE2fFQG/Cc6foerV5OJ2w3ELe0s7SzogCvgCOHrWWzXGmSskecFq8YtjdB7mqEtRekG
7FrKakHv9BswRcQDoa2HUMdEVjAeAuu2PMS+mSk0ESnlBEOsf+WIihsH0yEWZAguC5eOTqbu2ROf
o8ULzct2dCO/LUrc9OaiXZJesxroUYLKPVdAozftNakBq52b0wgDnXPkvV2lYfEyxG+EOwwxYcHC
UAHK+aZ0qNBxG3EGwdtsSyEa4t3sImgJLRxk4/eqdfvHGjjiB1v8bpttQSXa1NmBTlNmloclnZwA
MYuly4aVL9i3ljgx2mi6CREEXizQKLIzYv7g6z2NAjKr8tK+i75gWNFbOwYhefCUdzNKyWuQ+Etr
Pmne0UXGOmTWLkTPFp057g4gUZf5CACxl+hR5PKrhNauJPDcWCWdj0mS0wsMK/N2NtwkNPjLQ0iF
Tk3bv2BWkc+r+JnK95x/ybNjiOXMF7gxu7sS/p6KeIHjbJLE4Mu9kd9dnlWx7qCbDMUy8LGmoTkf
SA2tor0QQyscBy4nCkoNukE6JZTYK03GnEI7zGE9v6eUd5FFllsK+0G2C1Vt27Ug+/wN++fOMLnV
HSbOIkzl2fIxRmn8E+pRqk5dcOmXNUXZ5uq8Ea2UjNB2GHwo2zOHWn46g2SjcrAH7OoPy9WE6w4u
QV37JMwKZ5KQgeUiX68uK7fQDeAjvxXwf8V+tGFdBYxIPArJKHBrvedE8D/tb/UcwuxbvxdZQ5wP
9PhrTy6B6BgpoWxLjyovUdXnSS5OtGwWnhsFQg2MNHjlxbXo4ljoEPSvgRSNyVFMzFBqiEm5J4CA
W0dLfukvJqlXY08QhoziRGZsvghigMtLSuWByZ8UpUifuaFcF+8VYNTNP3ONHPVrKV4AQoXA6WbB
0RYi7FyDmrgLEV2Fg0SSrwV58rv0Ay5ae46UeSQdQ8qP+aVp5KToc4EX6+K3EMqxwGeJTKElGskL
YDe2hem6l74vHUoDl+l9hpn62jt90tJy6Or0nyksJlglCgFHezZ6rXNS8bdVO1Wbq8yLdcUYOLIo
7IJdvSel1jkETfRzXiKs6RUVQ5PzRrHbq/U3SP7nkDwy9wKmlUeubRL0WZ2XbP3agNFO5RsvltRf
Csj6c0fSl8iXEFC7cKY07Q9Lh5EcOO4DlThA3qPt62i7/2Cvz9LRDSJpClfE2xTWhhUVmv9Ry9A2
xPkW+K2p6FedldGPKgFdYrshxg76Kft4OUok3cl0Sji3ZnKtt8Pk2XF2RYqj8zJaBKE9V360gkd3
FR5bQ39xkyqeL2NhHnucJ7scAm/p+2PX11MzpX3gsn9p34wQezwJHAaxSp8NrzhGUf9FQ0GvVaj4
DmEv+/ylJc0h3MHAIqlpBEb9tKcI0qw4h1NAZ6fvWWOK5/Tg26QhOAbBQ7xMVF9Kd2pfzv539ju4
yr5vkG48DKLI/Vg/lTZBT/Uy+j6wr0YGri+aUXalFppK2G2+f8Oxbrr04iLlC45f0vdQaHGxa+Dh
PkrAsIFMFZEszId7PiXUGjrkVd9pTkJnE9UZLxEaXfyOgilNISnG7tp7tSts92sRJqK9buxnAG77
/tc2o5LLjnFrzHVhZ6C391QdUz1MLRk6EatAv4xma5gs218MWerLhznnPdBheE8oC5NbgiyB4Dwb
MDpVjc+5iazlPuHrlWSZY49nC8Q5/sSnfkCHrPXcxYa7xfdh0cNkot3CUWAdgwI3TvBduJBC22nb
TuRj1At79bcSH55RCofrwitrC8P9jAWDMQKSNL1bgfJma6E6ZD4lccvArukNHO9GuonFVyqntNsV
h8x/4lS2se8SdXDpvhI2yPAP2AbAbkmXSOInLlcB4Pz72bwZmXa4w3SELY/qRP2xn4EY0+plQedi
MMaVk0X2ZBGTlOGz8PzZwE5zU+zvN+69arHb7SuyUn4sLHxArLpb4AZzyf4Wp5sX8LUUhDDNypA2
Boyg05PC/g9OMDLb5FtjdffSxGGh2QA+s8gNzDImHuuuyqlP6RM9mDdwjKRWXDdKSriCBQn2Lxsw
rbCAy77XHJdTPe72cIYBOkC1HJg/BzZTTkh/k4YNZNeLfoh1i9bq/Sq6m121BDyifo/7mg6uAXLX
tO3nQ9rCkzQqAgOVmFk52gM+a6XBpYlIUsYCLea3RGRfkcfQB8y44jNZax9TjBeejPidYXmjVuIu
vhYAeCHEujqxRNYXm3HQsv1bKwPs2Ry7Ffgw0Utg+mwjQsBi6nuZtP9iaVLUR8fc9WRVf4ceyQFo
0RimapNMToQtzR8dEZJ6O86qfTZzzp6CD58sanhg8W4yZDRJmvbX7UZ4JiktkufJlEt5zBX7FcbI
k1P0hAJ1pX6YvAk1DFRVtKBDcJT+f2v9d9mUpERKFhPPkeVdIEeQ3PF+rjycq2O5SuFa8p4o7gSt
ShS1VnuiTdsUYqAPf3NsjrN7dutDytOKZUu9vtQQRpcQofcV7V/gqldu20NPBq+j1R+JpM0cHskT
l6G+SYfDvvtBjnDDtuy59jaWFVqMWqqvKCKfDwbQPsXNti6zuDxoIaz4gDwPZ8eZBuCOL8eEE3yt
Rub9GgIgAvAlJ0AviPQ/qPgRxY7jp6WzxS4UFVwyFRc6AHW2kOjFPcnqiR8JCDUJESKGMmORJfrR
iJ/xtqEadqx+gxS5fnhju1YNGEUKCYj9OXIJcdioRUj36mKpPrwyVy5HPzyn/zilzXDZ0VJMHrfi
RrUzeet6BZ/R5zL7lMajJb4nyHcXCXjcCVYiXfb06chBOnI/xjNQgHhqhHfR44IEFeDDhAe6m+lF
kCHH+dOebLgOM2EpPVTzPPT/VgECbm7ZoONo1oqlibRl2zQcEYqdwV6RwMiZCM7dvZHENc/oNbIi
a+fIrkXLT2fPFaTyc5A2OVbioaQ/6uWN70qbbTmbqFqf43lTeUDmIwwrry2RtjBYYve8cv9YqYri
pEz6QhIfqDixRi6PZwsMHWnqDumMmlmcJUdJuewg/QaOxpTJ0PKaCM/P+yQBfEQkeUzqHfz9FG5Z
gsf6crnPcb0p3mG6siE5TxaORsFvAMfzV9reSugMc4WsYk/CLGh1cSZ80ndR6lCZx7pRb7TKgrzn
4yZKNGs1OFVuTEQEOphXz06rnmd1rqgCqLX8TrfJFZUFGGsx9H++nTH0UTWVT0hIQi0JCQo3J3nn
FwsESNnETbtEj2LduylX6OQCWvciOkVovqkgyu7uwVAkPnra/mPAeCiBf1q9Zq0i2WoyaUqKtOT9
vjvzplpmB8pUWwxpBSWx8BOPT4ddHZw8WWwtP8bQcHDXhl6rAoSatce0RhOcz3VlRYAU8nEXMRkd
sijXz+RAXfOC13O13fRAU6DkUmClr8vHCNMkG7Pp8GouR02REWka3Ny8ehtseEpHBiDIPXk+IqIl
wNhHBsARjoin1h5QB9YFWRxsSneIGpk1pKim1JFhI42rNs647au9FDEuFJFNniX/wQW4LX+X7jX/
jEYN7t3YOUUF/Y6T17sXOf8XKyzzCCKFDvRRku0G8fKkpf8zFiMBsnGDbPpHCz0gVkhaSOAF8zy6
VQQkzWFsd58UhJ/l1+3xxN7D6eEsiLl9PTt1Vyor5M3Ts3lD6UNz27gcaEj38+0Hb+4gCPq3tIeb
EPGK/KJClRlZZDM83mvtZqmHo9Wofcm3IT9z1UY2DDI+kLl04ta4kGBSbkMVf05tkGA2geUYxxwO
ivgKw1X2P21PIOETZDVZClzQhuecaCTZIoj5+2sKOKvHrdI66h5YbNnr7pAHXy/EIveWxU2sYB0A
DIsdqHl2amKgNqYaJjl63ha17j8394d5hjsdFZycTK5m2sYfEOUIez71lNuWe5bAd0lqvpjwHyMc
gm9UvLF8amrDCb9BsCY1Vo/C0hT2WzlWt/Ck1VDoUwvMZ9ohEoDWYznfNAzN6Yn3Qi2DTjVK7QiX
ryTPAVY/6dyt6C9XFBapMkb5qnF58LxIRlqKNwCOUxRcoPD2K0PE7y0dJl4A5wP3tRLd6aMiP5b6
QrJAeiCoMEPf51Zw7/hK/Y8vcJZua1aOndpwUVzFLPkL7FvIIckkfYhzZYuVHU/9rku2FhAZ4dIP
seJGUJnsxFUby+IBj/J8gyEaZB9W+b/cVE70xjuey6CKbHg+Ha7EgMP7+j79guY6scSNN0vTgrxu
5I+0U5+johMtEJilNLIzhBn9pR6AhLisIp/QU9LyEEOLUU+onZON2nEQdc4WLv2dfGE4TJqz+rER
ptSHPOsFTm/n3eUu/pdpZoNx29J8+V/vOiG0W3wHC0a/mbvm36eHVz0m57vu21/qQ1XGtvlcl4RB
pKO25lg1qXlhVAvkGSwVAaXS2XTXlDjIziYqYVzx6BZCYIZNdw8636HNUj3racBvtXld9tG98dfF
kJ+Kb5iV7SvVFUlADx1GWoDEKrbcT6gSUIwGj81bHrm8I4xptn5+rbLD+y7rAYLR2os0F0KxWOGt
vweMjbyQyrXmPNbR0WlupiF9IqOzVTsbfkoYrRarwT5XtdlieD01QAeKERZ7GL26uhv4/jTwFhgH
rxmNldpnzy3sT08waLcamO+5K0mc8J6W483qgd+l91L/IhndMKf55JhVxTtZURQPexVIUyqUleA5
b2eXqSo3Okf6UTYQBMr7cxT+rVgv1ypJgkyAdwF04ivJ/EKrckk3AEOP/D2qjSnMgJR2Y7hRzy3Z
2XSXnt/3/fOLSZmwSpUoSWpKJOwPzWywk4ZfITodr8csft3QHB8G960pAOQ1i/Pp5EspOup8TsRy
ARMR/GS8gbXcMecerhsT96T8+rKIsMi392FPawq2gz3LCcbglWpaFsIr+puf2j50giYrmsmoWCeE
oYJsYClVH8z31IYIRFCcZVVBLY6gaPkJEmLKt667nbsOts7UHsb8WsnCj48BBztZFLMu2JUA7FZB
rX3DYTXYmndthLTXXQbIMb4l7po0+FwVX43c11BYYk8xbhyt10/kGO+CIQYJYUL433WM9kkw3yYR
ZTwYm09/9n6iEkoC/ATrpIHi7g9HThdm9HgQeDsk6vg4AbfBGcScSYpkEXX/6FV+sqpGTAfqiYpy
kwOAScPbD9ruQWiUtHe0RmHDdWZSTVhLH9btFXYGaAdQ+7+cyrNqP8mc+ZJcmWg65gRpcIWrfYon
7oG97fZzKBNtXFJ+Ab2vFkfHA+TFivccrcXywlee0oPfVDZHfCvSOf4HQOXueBoDbAMabj5H6Qe5
BugWcVypLfi3R8B7dUqNOz87Np/wtBP8DGzPvlYCFY29qFWgtj5PVB8FA3hJFit4syL0sMyaYP1t
UjMC5QIIh2dDmX//Rjf+H6t5ScG3YADF0bfHwrPssLiqO11WEsvYDFiwwYd4l6UlyiGiIrsPX9Fi
R4xPjM1oLrF2oc6eAIqknE8wR+xeVirMsAuCYVdI6AlxM30oklkw2JTcaosd+2b+/HUnXJaQHxNS
05zDkG3R6+aFNn+dCHGc+A+KWDC6YxkZCyOML6pPbuptna4EYgTLTHdltuKEE1qH7bcBO4D7KGoS
uRBJmNfnCU4nChmihn6L2prGa3/Pht2UP01DjQUfToJ4QPVHALY5F4baHe5jP69E6HosVEzWxvVz
WO47qLg8L4WffmPfLPGpsZMNqd6VPVOI951U/o0gslYK08Xi9awpWcH0T1j8/RHbMU93FtQutzkZ
+C+8qVPp+YZovEd5iA12jjIdT4Rk1sDqzpDe1TU98PsFJAP5tMFC/YdZaBf02OFRdlWMpx1jraoT
SBmqCK0Et1cuYWmTlK0sqNdJVDpc2UYbuTrS4PrGEIXsV75QrZQkDGeAE/2QRJqFxXjelQyXH8DX
+R5VPgb8gWL1P+Uw/x6AJWwVMsVXdTq1AnIj0saDtSgsK1LefMsc+fOKdilk6Olll1nh5J13AxOj
vrN5SVOLarVHjPKQTodwle+JS/+lNIsr38viH3XK4x68IwdHCV4aeXlOvgdYQhxFssepE1gsXAvB
QHT170oxYRu7wIpTpwKjMoZlku4s+GuyGe8TOazn2InToE/GgF2RsANLezkntu77uq9hejLwZUDC
gPzKQABsApnyzOPEy+czC0Mz6i/6KV/D3ph+Li50v2tS3Ogu3sV5f/P8aWvRWopWUHW/gCJFqkso
UO7ziUkcjCZu4SYmBkHRvv2CQuJ/ddV9KYQqkJ1dLXqPOjENtfKsMGaj34fAxe+SdmrI59tAfa4F
QJ15hHTd20AoAMcylDN9FwHSZDfsMUc1BZSCTw9GJvab23qVbNCKOdNQ8tnPyEKo6whnhmdW+lma
mWxCe1/hIAHuQp8W25uzkfPL39JOR55eK8lc8G65hPx3eLppcQ82hMu4Rtes5RCavfC3LO2OM87I
/26d1Td6G3xZJpGlIxe19bNkA5JmZPVQ91O/T+zsKH04Oe+ktVlSh/+m2qFLMR35sEdDaGU+fdwj
H6wLfiOyT6flmaR3hjZSocSWlOkISQB2qp4EIYXAoeCBsphJFqSqWsE5flvm/r+kaG54h5I2NuZD
Wm3geJqzEUAw/DbvJrblJK2swqgCIS3QYx3CK/UgnWa+047HVsvdZnp3kYWzyhQAMoz0eltiMFKL
QtoMyG4/JoEapqtN6Ee0Q/mMF1lbitQpf8ZLj7mE5MDskb0wY48rbP/FNUAMzG8cnhVrVGNP56kD
p0nBgcb5ixZEHvzlPZy04UXcndvJUh5y5fRpqEHHXCwRm3SVWnkvI9imNXSXdF319plQXPYJeFkv
wVit3O3OAlCttWpiQ1ocw6xk10OF6F0+dBlV6737XX8QJKXpB8JuTGDd9tLqG6cNsfYm0FkRHvTl
ZSD/WuKBFB5ji/F8ahy7MFZSKV6Gs9MLQlYysRrwUi93OzRFvxGqZF8ALxSqIfhcz3Ik5NAZUUSJ
HxWQCUY9IdN8rmyaBAjNnxTPPUoInn8h7QD+ISTXmxiEktjB3dwaX7gldHL9DEHng6NBQGAaoCOx
db0Z0CnSJKCIa8SpAsgfosCLLnU9my8ZfBynBkQAigx2h+RrgNsghF209bfQjDhBwT3tTmwzCxog
+JgZLXjTGhXttvpZapiUCuIHzG9hwqU0S1SlZcNgK1n3G8x4j0u1lly1eC/jceQ0/7Rc//NtyWMU
kw9E0N/aJB5x5QUsGXQqcLIPzD6OYBzwWhH1qc8FxR1BtgPOwwv3upQMvrbzKY0VbkARsjBiehts
YhcHcxHTU7Ew6WkMiRqJVyuuYy4RuFwCLkffpiAwoFsSLNvkP2rJs0X5c8mGSVZvmS88Zyk7usUD
NVeQNTk7aTzWeLSCfkYloCBuASyEyfHIbY1BKkuBmvj1KspAcje3PFdVRGjcgeWNDAnkGDD5TM4S
PsYuFmZTICqIRbYaiE1j3mV/fY0rlAfFEF/Si+6RvocEvjbPVhGe9betVEVt84S9v4lBpYe2Gh7J
a5bRvVwRLAJMgzt0euUaUn1C9sqPtsTPGnhsowJMGJf/I2ydCTdMgum2DFEt8KHIYQmVx3LiERwO
xTrYkwgR/0b7rK3zKNLfoRKDc+PVDAFYSScB00I8hamDfsVqk/vDTXdFKbqdg94Eb+vba/JDLjB4
XYWLUx6IEkRE6M5rQ9sgJSAdrt3NEfTBrW1sGoPx0lOG/Mm1FQrx7bwL5AubwVaRYvghbxs+IzFu
jARgIF3xp8Tgr5x4B6MA72nmMmuFOa9ro2IEpyVE/iz/VM2iSkhPeEw533aBJz0t/H4j31dFC+1S
gLOMNU2cGaQoaob7+vWbW2z3Rkbd78pyQj9bjXdT683Gt8nS3DREs+TEEozs5UR+QOHN7TmjNH4W
2PPmaRqvl08SxLNAojETN4ome67fpyH3XfqcnIhdBhNba3navJptAlScABcKYRrF1Tu0ii7iNjDN
hCQhL2+Pa3zqgh5UMXi28FOivtfsPFiOgFlYr3Rp5s8SA35gwsCu57NyPPWIwSb4unFk/lbt8iWY
afdzMbvgTjDF1wWwSBmLAZt5UwPbSGRZlYUmmBmeecYhv+AV4J4yiOGO9r82tQz26Kg/XbVkHO6S
jqB/L+7dOBaa8v+Kt/RTYuoULhdiQQAutY4I4Z026NQGQUpDIOFQEkoFcBQbAaHyUcqgJjXswMfY
Fmcxwytha/BPR2EakATtEEgA5iy6imqxTjjUeru7UpB8u9fku8YycV0yPaLMDdtkmvXmgxSl2/IS
jPlIGGifk8suaHoQ7su6pDqiOZmj3nklu6Z/WNPYiCTWZH3XQVh73C8oma1aqxXTAPaKLvGKPTtM
OefbOs84zc7iP7D1yXWhwerSEUvwfqqMfY9B04SplK3T2RdGc+OQBTVNaYDGBUlcxGSfG7Cr71Px
rZtx4T4DeYwtiNw47vr8juEGLlW9lhJ7xiyq9GU/K2ModSQVEZ8/Erc0bGrVl5xRlHXoDCfn3L+2
qJTrHIpOzChQCJSgcHJDovYvzMjRH841SpFswQsosddHspcX8Py2Huqf6sxOiUhiOZspl75A+068
tZbkOjNZmY0luQOJHAY/jVpL4WX0m5EHod38PvafKrop7iez4hH7Vr5dQ+kUjdITPvVBJ+ei1MZR
oNeUKQa/gH0jGhSdj3HncijlbaPJvhh3p4m9tWB3Q54oY4T1YINpBlfqika+/H5j4d1oliP8YE2W
q7NpeEpHjEIiR0Cnj5jvB8RJus5JAS/5MDM9wgV9YeaLijhx+68gl8BWSv0YesRX/SMkvaPoi8cA
Wdau+BUUNP495o5ZldoVoj5cbMANl/1N3ZWIEodoYgpFOEw1AGI1dWLJ5xqa87sq/iybGDeL7FTi
8jjAMI62l5pNQXUrZzcHCX1l2dHS6HfgOW4lds9alYP/++tDNtq+ngYS258NF4ogZrbaIC9pNXuY
P0bK6alSY6AJKou8Um3uvM4Q5vhuFtTDWZaHtTQzQYAXH4dRCnx/GCiYLyZrq6m2paD2QoLerjFo
9wvQ6LyHPS3oIi3Vim/Ua1qqEO2nREsU6E0nrJc7pV6DCqw9RagCtQXoqIngCR0YgkhGFJfpeEcc
hppoL/Dr0fIloPigjxQOqoSax3MWgL6pl6Gs6/+QK1relHiNl8woRFDPvx+yBtOnz+2cEtMOEEyv
L1qGJrgMF2h+ZQPLsMamxPVtE1MPbtvCigZo9YITMr5HU3eaiDh3FaGHzpeY44xXbpMJt3sJ5+SN
rAjoS4+416vr/5JLw6nqrrRQuhDzZqAAjyqlJikFG+zSge0YY8KqUqTymmHktqm8N40s6t72OJ/k
DZNbtzDrod9NxJwn+Q1PlW8jw/wCnr3xLjykYu9jjoU9wg5hwiFX4IlbOarYdwDVsoUyrSJZvWHZ
0JfXB0akrBKW6j/WF3V6uc3U8e8r66oYQW40QgTWXDGrdPHeVEgmkse3Cl0UqFvKBD8XIHGLeNQa
lvn1IUn7TIHwTdqSJN+PdOKb4l/pz6Ioe4T0HecscN+5QyMDdgHeD0xAbnIl1QRrYyGCQOO14KZG
5u100bjKD4oOTU30NbLnpFI+TTlveqLxRjmrz0yu5/CVIZpaWJo9Fsg4Sspxkq8bTyH29hRXEl/B
q8c6XkYiyT0pKIitHYd4LNSM2pO9ZfhXDLLADt7SSLdKfH4oLtVagYbPIO5OSCjYOEYlfkBvuxVT
pA8LtJY0nGVNiCoqADBWh7LqfsGKF4nvXN/gZhGudEqupJfCAr4xCJNitJSMHpFGFDcEk9BIquDV
J8Uan5dP2OUSdxnr0DJS/CcadMPR667FEGILZuD6m6UbxM9f+nNn6w79f61MSUi/32CHPAvxdtr6
ybGmDOKm/pElDYV+DZFNv4AYL4xA4vEhrFYG4ci0ZWQeSyynjbfsQUc6U6Qbn40bng38+iG7PYZj
r5pxfVlh+kS4Fq+3uvNb1mIqvARBtL3oKsInfYSM6PyU3Lvl1esLPy2jQchddzj6HoJWmjZg/kS8
sQg6e6tt5q6XKzRAOVY8NTU1Vngtn0Sl2tjUumdyh8Fly9+h/n/dH5zSMUOBcJYxrxVCcoWlidTs
fmAlUM5bdTFG4SXI86m8w6aXt6cEizQznskdgN+h1Vc/uoAAOrYgeLoRHSrYetwwL8qL+2ScnoBm
W/EYa4Mt5LyarIpIyAMZIq3kToFzjoQhr0o7pCUFb+Df2lXsBMee0hRj9I0jDcKbxmJIzI33erWT
PshXXM/PRm2IHG6e+Yu9ext1Y4ucVqMJKE+CnY5uoG+p2QsD4SFlWJfBb5yChWXk8uQgB2hUc0lH
sk+82XJ00ox5ZG9zSKSzn9L8MFMGu1K5v+WvgMz5e+eGQvdtbUloxnQEUkQ3sHdZQdqwgsboj4Pv
JHhWR41HU5yu0NhpUfAyDAjEDK2gzwVfWCWziz72nkG8qPgvWT1j7mGkCzP+6cZHW0driRobVweW
cl6DzZcHBVpyIXwvTBKouUIKDRsLureSKQgleXlEt3YJkQkmbyG/oaeJeMHOPZSTW0UkOxeZLnft
YcHxpPoE6ppM06o9I1KnpeUdkSIDCQk2YiGWC2k62za4Jye99gJhNv+Z/4WRP+SZMVoR5mJw+lY9
L9DUs1AnjGPFBBBuXgMv6BVQdWbOB/xkS/lbIi625uC0cU1LEGh3mlhmT9++mxxjTW8ht3rn67H/
/V8lpMs9Cu83/i+jO/ojYOcwvwVygTuiygpzHgtm0rO8YCDqnqevNEP8ZvyNWv8cib6j46wUvhpw
IQivy39C4tH1TdqM5JDV6E2JojEoYdN9pL6OoE1zYJTIiDxwflWasAKLS2P8JpbgGxDVV1JIS5N7
eBewDyvxH6KLZEx6Qh7rG6dpJGolq+bv9ofbGtshDTyIuOD++8tj+SIfJkgxr3dGLi6xDhCwizbb
qGZUH1snOHW4LWtgpaMAaB9cCEB0gJe95nEbmw3ldqZ430N8eH89cbfzwncFz+BJXu7t7bJUlbk5
LG6rXHUd2ubLu4Y1+cZ8IVqCP6QEWwDeS/4tA5EFlTxRVmSY93LUZEmFn1r+B1DBAb0hT3zSVgbG
/VJzo2KMTZF+MYAdlDhZwr/vxLf0jLKAcLMG0nye8OjOFP4vSltxft5uZouXZMpplC6+XX7otpVu
F7IPlNQmCYN1Iz0i4fuRuX5sR75Akmuzf5+ISr60tc1PJLQKYXdjXT0kJLmKRAn8MPW379azZ/62
VLX7VOSzFbFBOjlr0IAz2syjvzYW+m3mR+Uma+gMngI4kqVYnWXE4YAnARzjiYv1SkayPtvJl9k5
1ISVqwWujns6t9n5XDahFRBc/NJdOGnsEEHDHFt88wZT+1OVgRe2OefevLUoZSN3sgY2spQrn6GK
n0Tts73p+fEfu38yujE9O+Mb0DxTjhp4kJsD/OyDw9VFhaz4V/vophZww+hctRlh7oEEq1HCE08Y
kgr+zMCbDJou+oqe8fsvj6ulxgT6/ClYOzGFtx143iTIVQ4IxS6iUkpU1LEpltzJevYOlADwJF7F
pj4/reJxROKVoXfJwJvLbF+CjmCr3xwGs5gxKdgxd/F5Lpd4/t9fyEiHmk0WyfJ7tp5l2xa3KHyM
VgiefW+7/ZHgUFu21cINnku7tkAUyDn9cVv/kg+c57cjMexYbqjBRHNtmQS6jarZj6EgBdJHVlxu
Ge3oDBu38N+6UVFN0vNeFxKG2y3diLj83NgvhbSkunNgjanmpMYDt6cPCX+g9MApvUPHoz9ottmx
XXSG1wmZw4wGoBzO+sFGc1AfGqfQmvDsOrFaSgPC2jIXlJVDly2Dd8fVm9UdtR7lkk29bauFuqGO
qSw1hdq0AJ40sxYcQsG+m2uK4ZeElTlhbu856McD3yY5qJNTZZOQ0uzV+nIsTqcbmI3q2NUB3bxo
1daWpHWDfNdBMac5JukTl0WQvwk7bsnLMFtE13KtpIcAmN5fTtEx0Ha8vavJhfsbh5ftGl0gYhMt
oaN8fKaBaTsbf2jhDn9R1ml/daRCg/Mo7GfXDidiAwOOSA2lOw9ClEYTvGCnNXGJvJhOr+4Io+dP
gyoYL7A0YapF5e/xux+BQSAXXpBUwvE6/g+JcU8XaMKJhJBabfdhrmzND7ZVW1viUf7r8oFETxOH
89rPH45U/VMAW5MdOdq8y2JudMGCrsrlz6DEhFO1P9Z/2LTGunfzgQJGNaGzTA6PfK5wx/Ez+2Nf
Mn4ohqxPI8PCj0acyiq0D3uCKZ85JrP/g3s0tJvQvwpvaQJ6vvnbQXvvuIQS9h2RWdigiSfJVTfP
OYDlyvaktzsfBaYg0aHAzBSEj5hKoLL96vQ72Ll1Zo42V+csfPpvpiMSLhFt6yeY3vY93q5e6ZLd
QWSA0d2yPe2YNT1tnY+g/JyucsyarsmEpmcqjyKcpF2szolJNQOJSsl99pOwA9/KNjmYU2dYj0Im
v/q6aI1hZw14UhhLDi5BaSOJVKIn4aLVUSk6oRybg0+s331ejUC7oCslcJEUMIQM3P2ye7ChFCic
I+PuI4alFYjQ7saHle83EdAXmfsicCW4tCxY+odoDpXFYIE2pXgDCMERpLwKA7JaOImQYhIInAOb
/HHd0QfaSca1Yvnra993FkmxrsuwbRVX6xq9OMAjMth5lyhzQqR2psCqtdcb0gG9PN51l99RI9/e
l+oJc7hXPmuKORdlSsMseggafVN3fWH37VIkO7W+N4c6Cr8XGEburi1TKLnEefKsLl2V4JiQR8sL
FuZ3Q7f+70XwvaF0Fj+qAiwHPVWY3LkN00CSLUjTqbER7aTlv9ScHq6f3QDj/7zwJfj7hUIU1EUU
2fZctDRZXpvPljYBUDGz2rP/FR6HmJK3dJ/9+AfeHWIa+jxXZo/N3SnGypdEs5rKM4SYQ3HNfd5j
oDwJiix1iglGOVSByHbkiHo+7n4p/moGtMPL/3/Psti4nY40oGZx0gB78HP/HO/3UYnD3SZSH9pW
SE8zHHSB1aT9zzFIGrPG7Bq4dSDCKreC1rT+p4sG8+wQQ3BlNiM3BWjbfjqkeyQCnzLVujEpD63B
SQocEonFB9PoqEHGdVYqgC/kJSvVDqekE3TTV9jGeXZKN9yTRO/5OaTrKXCqqBk68DWgdzdAuANM
kcr7e6Tiqz1pLMGmhKTBHLYOl8FXe3EP6A5ZiqDJWjTmhzIBcRjLmpgAqXmKFV9klXPyEMnQW4e4
OhVJLcAdufBaKyNEUwup3ECVTXjl6GMkR9xb08QWc1U2tK1AkQlqyu2Uw6QSyfao1cEOd8SWsgbU
TVeBcPNu2vDXIkeHpIqXjM8Y5byYGVI9VPPDEupU2OMmxPyIitrddltx4WuDcTG1F0PoFYp054JN
E/Yu7hXQA9Zd+9zxD2HIBddRFXKr9ahVheLJA/J/QOHYwfGXo8YfYYgNSI4GyT6bHkP7P6s8jEbN
COjYzIyHP5jc9Bj4JpFVfbY6pB9MtiZv5eKwSIkZxwLjkxnTregYfTl4t1BBkZJNyGL1YKuqAMeq
isifst9Ita+34gl9gObDj+ZHHqWql2WA7HNDNpk1taPMqj/dlLgjl7gNtMId6/PTnIB0eg//Zomw
av4M9q/zcviBvcKeXij6UDONpcfoqt+l/iY+us+BR8LY2yRw/X3pg8I7MS+ldqtEZeR+6c4WAO13
/dcYk7dFJTq1EAi2zIoxEtNt6iuN25UAxrS84xItNHkDlvESl6+Udo9WSxLZigMo4fztrT3VJWxD
py3Ku1d46SdIrUv5lGg9Q0FMSjHd5Kwl/QDdjpClh2PdNbwdaIDyJ5kI6vATKAx+CUsg5w1ih/na
c5HLvafc12GwKHeMUZjhQs6otuIjgL8TNkqQUEmNX0nVTd1+A5d64jAYeFTLC3VukBlVykN7SHh0
jkiYJx0NI/ekAqS2IjfF4zpL1WusGpGQSDjq4neRf0xG+DNsbnWzlE+4LxSRX7MPKE/9R0hpK8B8
YMlwK8xDwCZTWLdCDeIYxDEPEVLqxqYxkXm25uifuSeWug6offFsubUqUqNQxf//uIxsWseMphRs
8PIkytMzbiOM1aJ6ux0gQATUwWH9QdwMV12WlthrN4dJdE8F1G+UfQyIQLBBECjabEC35J3PqOk6
40rIHsEJeDWhgjmzwxKcZVS5vePhaYhASdwauCfRmpinCn8TlsX1BybNxvOovN7s/T7OtatuKHpQ
b4N81+7UBAt71cTa0fRa6U1LArzcLzQqgnsQmtrPRmmatMB0OwHVxOW8O5dqp4G4x7SSnqGUGXs0
v0dPzom0zXwJfA5Fe2G5MyWCwnLTGqxPqaMx9VSCYvohyqlFeXPJ1Td5USxWCZHm8+U7Dpm089TD
+4J8tF0xzoA+Ax7SMi9FRTM4+KSuTzSxQuqNaiiPo9Bef5oVIPP6ybhX2iQWAF8XywJtV2ZCp3x8
FAOncr0+jMS57GRjykMINC9WW2rh76lM3ylo5S5aVYP/EEcuzlir/EMyAu91NbiZIuV4JATy+0DL
in5neJwVL1v2rBDvUwIOMpSMY7Mnh3m64165a6eVp3udeLi4dsfdwZh6WAduQynarSXNtHKay03Y
uyE2bHfDbXXTgptW83r36Z04oHzSd4XzLH17AEebsCYsx36qQbnSrHObMs+8NqwXaVkzACoA2KEB
Y72XvphuS71facCLkmOhyHyC3WBp1mP4HV2GCC4VN4V8pcumATXjDGC3aZb3QIqf4Txix6HpvSWN
UzvA01m7E6VvyJHsVjsXMX2+V8zZXUS1gV6CjNhL2gtn3m3OpBOx7+JxVNXwVndDpcO0UmEIiT3N
VhPzmy70cWUoFZIEOVpeJGedxf/ZWzmf7o7LUjS4ZlK68sN9PGQ8S2y17eE7CGFEwU1q/wom8nLP
SB5U6d9MLDrZW9gd840SrQxdCRTd6Pm75vZ2UrsvH9whkHUqn9XtT3EiFj7lRelihy2a1d71eoEs
Od8LvEG8lZ8PRdgh7kvYV2v3nZNIuAKKFrXpI/rPutIRv7g9TTRreF5snQIRHSMb760eYZSQGK9M
OamSt1OGwlS0LHjw7atDT+/VLZjWpZZG8rDeDlk7+gHHk8rxmivFGh3GCfkNZsE1BRddn5RW24j3
tGMkmHYG8sQToqrXzQuI/JINCXGzQEjQywfDkPmL3HrfXkXqML5HGD3LBof7PDnOZgZ/g7XgIONI
vvk5OhjyOUqQbv1lZ/2i3k4tt7rY6scndA2HR4HqxpB/KapL+7GDAvEFuhTBHsX16ao7p/ADRL3x
zdI00K1S3TQNXnOKzAKeQ8IeefKUfXZwySX91B8TgXT/nN5REjcOs+4BkIQWAJAayHdA0Zn9QKMX
QkfXwrfI1/eJcEVHzGtgMj+3+AAB5odqSdWSPc2gKWZetKr3fVBJ24T50DnTsQWCBhnbm/pKaxMR
FWMjN8fL5vnbqAi9OhtNWW6OJfj5sZq/wuCqNr43m/kQ2pcaDDSCe2pLCnnxXRPvYW7qEAAm155v
GqgnouB2ONCV58QHQQ+nESnuGdBEMBGDg57AF152GgAnPd1wX0t3qx6W+rQkdd8heYCq5iFL923p
Gz8SkgwZEgaL4G+KmuRsqDhd6LXyB6h/l4yyYUqTVY9DfeXCMy7FU8kUtU2jjnuqQ/QtpZj3GEPF
kWTqKyzDtb73imi0XFwIXngWr3Tpc2WYo45rjM/F3MUewjSkBhNiYXiRSrVxHowthufPz/nwEYOc
Z4lENY4JMRtmQEqYo+e0akUAf1NuLOGtKeQ8wEl108LfWp32GkVV7EGXzC4JT/VbF6gZSRiw0dK8
4X6yVzzL9HdRMJ4wKgnfODjogTHzDZfBF4JAlrk3MU/2SnCa+DBiBuoLEeYokwrH+RL7oEfcyGG1
VuwOnJYW6aqXsMKzVgYAIzaUZ9Js3SPsfvRB14fGCgB59tvpoI3QocTP3wEbj/T0agy+N0M2kIp4
bC4vv63zAiCVhmGhiTIePw7IiSih6MX0HAnIeEluoUfnCpWSMizroSX50sh8fTSrcpjnwadDH+kY
4dGfU3ZW1rHZqK9tTfgWXKZ0fLji4Nj38C+jcN9idfL1YGxk2v6X7ZiN5K0JXe640rSBKUyuR7EL
zHHdCckv9b3l17CsxIJWvmZVtEH1tHYqIhxdgYsliegQDKulLdu6T5UpOf/RIG14FMn3zMA3gncy
sGugoeAuqL5ZGCfuDOzW+na7HxMEKYIYLQV7JXPpF5uWYdURFK4Mrh3IQRdqlb2GdEQljyfPLELW
E2Ez+7azl/bZJCB5Mr4uwADQrIgQqZBbsRQfwkegJ4ZtmKCPvLagVVzSwgWBdK25+ix7lD81PpEN
pOY3i71KcH7oiUQA2Pm1NARYH4uxuT9vKuuK5Akyyb80FGqmOjUlZxR0XbSkqXqk83AaL7QOFCJt
dFfH5wBB5fuuttVHF9mtYn1ZXAeDW43lZkYHzQ0VX1VAjQaWbih5i/s/v8GVDM92kOE9u8EHgDGy
KaH1LSNPA9K3LRY2Dwqn8/a82oEMnxSaOyn8YC/maQ2vcty2JgQTXH5WcHjLMXkIlBTuxnoaRYqR
aoBes+jumgQk8pbwiAuitBVQYRpZ76JEsuYJBvvyoEVnb0zZBDRM8YEKAxn8DhwNMjAuKgqX0hC5
p4KhVcbtqjhIA31scAuQLrE8/q3REBfbrc0YHdzfHuL5iGCoHf4sXirRdoujSJVEo0Ke00L9cIcZ
EcDnBWYbfJKD5orMKOPR5Djr6/rTTepVqlXtXaYMABWSo49AsLSVcd3wXHHnh8/i3sc9j2a4CWZQ
7oq+FIas3zrQEsaHgj4vkdthK7JMvdH9+FSlwoJdnS0+2xIoVS2RvqiTSETAZqb71/cyx2RcZin5
gulbvExFjom7MsXDeaCCnQCneRcNvZyjniWJ72y135IEN/i0xtpqEnm8pWIjimha27l6OTT+o7Jp
tEFT0dsCfTcnOT/PwReRiu7GF3rs12GX7O2DYupOu71oF8L0epZ1GACTd71UtiidxKZJpz4f2lKh
3snII3xQeJOWva/uOWgzx3vcbpyJTX5WfRmvqeLFJPZbaUPRcgcyMujKsfsGxIXoGQfoLlKt/tPA
efIMkbRNXd1EdAL3BXld/sJzseXSuWMiVS636A0dVYUSmUMnMR9EFNWXdRda9lpr3qnfc9or8VE/
KvRJpkSQPUW8xJLTSkQGAIe2nWMlYgYnyRGwAWDitPFpqRuocn2luRtCzTupRCQXcO50YUwxrn/y
axygGqyUhXUAluZw+8yknSAA3wfNoambVqBvp4KLM2/aK49V9s3f6sQz6Sg8W1/UZY3sltYi5fuy
9W6WtmDpZ2QzwGr9utCgP1aZTtRv+UQYQtwcNVKmVCXYTshY7EBmdNbYs4zKqNyd3FiReGKekvFO
fu4/GdmV/Cas1b93TGwQVAKuyKMVLCekyyuxmv3OK/cvQ5GbMwipyqTkDt61RxB8XamuZuEKHJNE
BqouTZlAIL1y4YvMo05hHcrk1aVC6HeTJ7RO01EKyM7Tmb/S8SfuSpQRuGAsfD4WXaSS1Ijb/0oM
oVM+MBKYZC6OIXMYWF/xncGVXbUF65j/ISGnNn2rAE290rFUvz2Ibjx/nfRzgowpyaZYj72WboVF
SP6KZiBlcjsZ438Q70btbkGYd6hrSIafFpMNaa99W/na4ojVXBWRK2NKhZ79YdgfHvllZxfnfANj
WVq2IcHNKTYGHXmJYhXg6EP2g2AvGyauJPN95I9/HIgoUbl3XmC9W3jQdkrF/+nwmZr1YbjA0ZlO
0uUGA1kBYX4xka+DSModHVPQ4vUN871IrwDEI/DJN1J08KH+Igu1T63xX70fjKdDYRkTlfIkkgdO
k3cvF0NArcY2ssKk6Xe6OyekAJtC2+SIYfjp8U4KldctT4J3MfJVfXqel9zB5dbP/evL/wNnGJZ2
lLbW/+7NShAVY6EVnYKHEp9EoQUUU9+aWXAoE8tt2nOl/eXKPA3HGAs9SqN+D7EfWJ6RqpgWGnOb
dQb9gqriBCBg9/sqPhcgFz8RkHcahJAngn/b8RlA+q6BC9Ou+8sp3nTk62Btldyk0ffgPmUPs0+G
EUGFWrPsL0omdLwWQlhJPOJY+dhHCc43HzIiIhnwoUyvApaCBjmZdEyB3hZIkSGoIpdTlNDx2lRs
ivUHKyT62S9GtueGZY/wdqlpn1mT2lD68j4iQ9+CsLCAhXq/GT2XUdzqeg3o3RqZSj5uuIUWrN84
2Hw41ZvkGjlfbOmjWEnejQ+RA0nqjZ8L6uS7SbUUaFRGSFUuWdxfhza0wnGhdomVUmHK+fD6gC/H
1SbQ/qQ7H9+VksvlRdtAP+jpsF9A1XYNa7Ys7vkfpyxaRP72CfbnjWTQCbymRHh/JjSiQsLhwF/F
ZTfTIZsfMy2T/35/k/vFzzjq6AWfR3dmPgCX8FLacEgUgZ7iW6NWaCFYKz7ZHiNnw9gmNalTYE4d
1NhQR0jZ976ItC2E+NW5PTAubdYIZTy0S5gIl5ZyqWGSzkIjGPUlTmKbpJB5b6OiXOekBEzqhOrS
GbDuRVOBF3RC+QaAnclwg6ujbTh5JYsK1B9bI1TVGDRkGa8Rrde4tKSVoOaVOPqcLGjUCsH0sWWG
lFOb2xqYYhQ2oc3ajcFii1gFUsdmP5YsB+A3VoaR0XTmBIS+ePhcD/x+a4CFvznUs8aa450zeXWt
3mUla5qZP37IRydhNdlfrCoXJH6Rl4/omm5twjNjNWNXPiAbKWVsHdNdNXKXFSYnzR0NS4gZAIXd
/L+I7zRkm/SeOGyXxQMuINAmQsZRz+5KeRSqJBs7Phe4HemartPv3ovGghpn6na3MaYFUN1gs5sP
Ms+VJ5VQrJOsNKFy+wI1lfSLuh4CXl5HNiarzVxnFwXnE6oB0xmzhOGPGxXc2bXSsngFzVP4HEzW
OrBvv1PA0y3mjEMgIhA3HZ6QkpRwpyCNYthnUlTduS0i/UARM9Y8w+R0Nabji90mhMS6TBgiQ16l
wgeZvTD+Tt5wQxwmkimtkdi+IotzQSejVzD+xcPArh96gWfYDgXrhRAimxh7SWv80ca28UYmmQFQ
yWYp1NQC2hSvt46gevxIN54gDFV0TyWpiy9tFfdPQf3Dnyo5kTsP0AKfenHmyFShucde+dJjm2sI
xBTpodm3oKodE9rLCjt8WUVLEbAccd7+6JK4HY+upqup7L75kZQ+rs/Gf3KAzFDhPo1tFNT76tW/
iz8atQHjzLvrkNjmTKjucM1Dz+wpXLC1ZVmN1wYUAbrAEe5QwsZLl8bzdowsItcVmBsGtJfquU68
c+2K7F0wRi0BnjokwRBVzfhafPG/HnhtFjxYqCe1PNK/T1beMpLkyQ6cOF8CZfplq7XNxyuJxrTr
YlpS8SODF8JFjWO8GezOcNGfkU2leVNZKhdVS3YqcnQHtJJ0Z5Zf9EQlcKcMkDg9yiwhg/ba1iO9
RKQ8bUXaVBVnDgkLE7EB3igcYy/wpW3tG+dqg2jfKKSEhETVruxsBluCRJvRciFbahM4Garz8VXF
IV/QOrAXIhvVYQZaYdRx3hzuP7SzxXTgUSq48c58nJLxVUJFUW4IO40Ah0SVov/vdZzkZ3a/GCz/
2LnxASr1gY5jnNxZ8iEEoXr07muAXZ1SCmwQYDScZnoez4Jhpmeq2ukgwCBaQzj5q+o4VlulWGCQ
tFUOHozVT8mcPdSrwE9ep++5JjmE5HVaDeHzE38ORZEwDhW8CEWgHklZyXNDqtfHL/rr8fJ+NbpA
mJdWBd0E8sfjewYNSF0gXg/gfD1ac1Bl52WCwgj1RWqt2P3NNvlDGmSHeOCg2CdL3ROrTTsQfpJw
fMdOZGpEuRRnXs9Ba9h+p7mBl5ICnQ//FYXIweQB7R4krxHFL5boVj27xBBhAcFXnnrGpLC0Xke2
VxnSxy9Q8fHk9f7MjYOlHvpkSLX+j3g6zrtawEZanyRKe/fVAYSsCi8TkRq8rhFC2Q44CYLMT7so
CI1tItacQ1yUqJItX3B9LxCORTK0gagUh80XhW5cCxNCeno2Bko01klWo9Vl5kDBH7lFeOKLpu22
N/X9CI6xx1705Hjhchy3DhlERQnwav5g3c55Paj5K0LelmFSpsIYvKKmxMB6gKxFomcIXkKxtVD9
3df0f2HV91sxFkavH7JZJ+7CAGOPxgAcKdPDPmYkn0483XQmaXVFduC+UZUcVdiycdtJGqOqJm/1
F+SJm2lTS0W256B2hn3gDbZJOlGR3jnTbJrRcB88MueOwpGlVJ8oIOuVVia1Gc1sl9ReMzgoq7O2
5wB354jAGLP1hI6hhlGnDxttJghWCNZ/zdTuTiOyztEW1xgN0QMWOHPZKpZXGg86to2QfoBmqy/f
Ejwu4XjbSP4esmaoievN/0J8n9HbXO1CcZ8+CNw1JIakulXP+NuKKxZL6akfHsdPP+q1VqQ4HuvE
GmuLFKoSstXZos9XxG9Shtx8lkRU5bOxr3f9l7wc4zq0wNtoNHYopMztw7hgEB2r0vLXO3FggmfF
zusTmWJ2Sj6BAPTVuQNPgYsnL0IHFSpobzB5aihp6FJTOSAP8rEmxJv/Uwu2QCFlN+ff6rvSSRMi
wgk6SQwCqSnpmplr87WjH+BBg4T8ajsKbfP0JrGEBpkLkauCZty31iAbAyzQp6PWRnaukqDGnDIm
OyPDChEpTrBnozNbyIU8HFsC5BsSnyybUknbbevtmMMN51cT0FIpUvPoE8pxjreZO6FHA8tb9ABA
NnE4G5tzIG0H2AvPr+wooJ1qlOiZlmidAG8gWdffQ2aPddYPc9UTdleGPiZ7P+XbLfJnwNvgaYwZ
s3UD898OLbS4uR3CqMdrrEaZWpN4BQdawdEndAkX5NJsf1NxWmR37E9jLIHdldncXTE0g0INR1kM
lE6C8S8JU8ZGjKyj5dGe1QookA63EB7GiENHpQlQS+HMMxhZU90sGzfeoqZ9DeCrWrw5G7hbLOnW
QH/ScNNaoz4Z8wFNRPmwf7DD9CEbFjjrdKRcv7QU1Xs9S8iwyVsH7mtPuJwolyFVRWS0KUmasiv0
ni77FS6IEbODPk0m2l/SU+WnRO4o5IZnpNyy2C3CFuix24EzV42RjJ9x4SYGb9wFXKcDWXC8APiT
TSHb5s6oO4QVxyK4EV7fW/OUZSse9bqBr4lkrB2iTCxWDTygJhNYdqyRJukA5sxlP21ADgqOx02q
Ivicuogbi+wUl7r9fW/Z0o/7bWVC2N6piuY3OGM7y/SQjwCyKefyC7DN/2P9ITARG9SpzWALvANl
+SehfkZdnArKTM6bMrHHwAR81cZBPMvfKFTFaIBAGsIatXXpfdWmcuEJO2pi4ajhnGDXRvoUwA35
c+T42ZbzO6cSVMRMjKtyMAlUtoigs8CMV9Ppia6Y0YqrVliSESlcNquJN9ejCogEL4joid30Ec0L
/120S/u4SLED4LkHW7qQjJamkdTakuu459Hzcd3h1alWhXFC/XKcBDaDivCZqA8HxiwDWJu/fovz
PU/oT7epPtX/6R6wmb7jnpT+uwr78M8eOMPs8OMgyDPEjW1MpiAbkbTRC18hnYRD6v9QJJLYioxB
7S0uJ2FmA6VyP2z3it3iV0VfBoFUJj+ltbseWchp7OYCRJPLc0cS/g6MHkiiROqzFCWMetnKrY6f
IS4AokIyy68uIz3NHaEfpc6ShntowXeF5KugGrHVqqBkLzCVDqAnlqF9V1AYby68JKyzgibOLWGf
XoLvvB1A33KOz/zBsXm54wGCMj9BD/2p5i1sUVJEdi3Db6fxxXmQaEQ/BJuN/efDodvncNqCGSny
OAFlXA+P6MWo89qmGXbCc4262uj5ym9n9tfa7g6bhSL4Hx8u74JlCpkEnYL5TC4rTtRE+gjk5Xks
YfHzuA3ApMawlR9Hi7wbq8zPxmiDuAiWc4l8m8cgNCbWvCfmjgK/QKhjL43m0k7cNeyn6TYISGeE
+SRGk7/wB9NZhqQ7c+TDVEMVV7oGAfZ0uPfyNM6xYPafLEQMsQFSJ5jOqTb909RXn/BXrGLoliMF
XU9tUBI4POanqFIvCf9c55m3KFXaqkqbm1AgPFqCnkt1c171G71O+38zfNwdqI/RMhKRvKPYp8Uj
3vRK/jqMBxrL7h7R/3exbmPkP21M4+acqQHJV8CtnRttfjZ9gGdKyUV6htLACJ9vu32mxQY8VP4W
AqrVdeBsiZv2Qnwd94Be2p4ob1zi3lf+i5Y/t2zcebm1qUb//1JfgpDuwznyC8GT7SDiIhCLxYmq
9Tc9pxK8iInMK2HSf0jmZtuNNuriUwMIRxfB3fjC2KYoN5tch9rsBd9bTnuTOhu225lnALNHNk1h
bhb5l9o/Ohwf903tAjGRzrIC8XGd0uPa/3MZzYWSeGRCL2RGpwOlU8f9hcUOcVhZdHFUNVvN9KaM
Z5KUXJe5d27kYMEL5uhZin9VmrE3fviN6O9sftxatMf9Qs9sUTOU7jRtSLXHjw88P0vIGp1n/GEW
PsVTymkJlX8oXpXfbFXaImrvz20/AoI79/waYLtB2ae+nGxswiBKEJnZR73i5MIUyuVrlg9SEVBI
ju4Dqdyhta4OO6iMhPZvRJgH3EkyTH3D/6Yrsktp0PcYxnuQxlOZNSj8NPQnea+0v/8J1oWQOWIJ
0sfTPAlncUam186sQtE19xvkS1l1pH05TYDVWveOQGhG0EyWKMBUKvhCvLP3uASt3cy4uOPphv0K
9F10thf0kXi0I+uGb+AlLFbyjdv1/Qx6hiBmxBQqnYiKC/94V2MMS7L++p6aiD6FXtE+LSQE4iC6
EiQPDAat34Sd0ssyfMr7mFnhuGk1slSy0MeghOm7gAgg7rp9R+s3bLJhnFz4bTiQLlqMU7vie1uB
R6SmbFOfJokifMi6mdS8Ub0Wy98hjloGaCT39KMhA3Zr3OtqL8IaKkjyk6xUabLx7eHAUHeS1lBP
5pViRIdyGGaq7FNpIk9HEqJFkQZ5LazsG2mduC9qipkrftIkc2lNv+j7Xuf7X/zeXubgXGeaQUu1
7fpymjLvXo4OzhGSlZ/WhR6oF6Uk1zOF5U8ocxObgkfzZ4v+64rc5vkT4DtRxtuI3ALYEiqwfIlD
doflf0M56Zp3JSJIvYfAsfRQ0KQJauKIG2+YJxs7GDygOQzqifFr/0PAX5xQ/l+XkX0PGtl37g5/
kIfaxsF3Blpi7rvj5aXXjFwwpkvZgLZW39qNhlT5cctxhisBAlvHxs3PrBt87edbioEXZOU7Jb6i
xzv7sSuFe++tuiYNB4xQGv/PGUo3Gv0FDg2t1zCdrDLS5tjCIgMJf+KWdJLzR4I4APh0E9cej/4C
gpKb8KbXEEG4mkygLdZl1vGMLUKdSb2LgVJwCemoLm2ghGwXrX2kZ3caITnUQl/nmItDOkw89gR1
8aFhnzwXWTU3QDiTuApAV/kMDU3w/WINvt50IjlBo7/2aeC85mYbrTPpnD56DhU7Ja1ylJXYO1Ls
hsdtAKzBseY5TZUsrpZyEucclkURB3LUag33txg5FnRZIKkucODnF5LYib4Z/UvikmOe++YLM1j4
9pSsiWyM6lSe5BTpOFA+PihIrX8whyAYXM+2oratzEw+cgVaWEKQjb9QZUADYB/SywrTeMC1S6t8
OWU0wGAFPdhh4KD8Hqmvxi6/4vm0vcjxrMY12AZA3RCU56u+wc/XfX1/6qU697Mm+7rf3Tj8MiNR
UcqNItfbLM9w9qbP0MtL4iyYncpHWyPh6B42p8HLMSUHDZQ7WJfWU0f2QdgdOnMo9KWrvX8q9LmJ
lhgngFsXpGF0IPU3bvOq89PCiDLpWN4yfBfa0pFC37Fbtk058eQ9ouFrwSTb4dQ85+FntFLaTAlU
cFQhxRbO+cEfWWHK8akIza2qukMQ9F4jB/MrltxKMnUAuVLwueBHohbxfCreqGj6mJNb+4u1ubo5
ufVdWkh5832A/d7gkQpCC+PhHJu5E12cDwmfQKkE9o58mnBLdlHDmO/PfB1cGpJV7D4PIm4fWpkn
GbGWQwjbXQrW+Fah5IVkvx9wViN53Jcr8IeQ0IWquLuiMfTUcTsI7uZAITCuR/ERaWnHmM0V6qgw
LVCzIOA9TSl8pagKpHLjD7WQPnJktGrWKSr0fVcSgaeBIMlSEGoilqilW3+e+7vVG77CdITN448k
Wsbb0vzOUGtC61eNA5NPrl+V1+PO7G5dD/AvS1IZhEmFPyC5NJSz81xSU5j15KNOW5W3GP2dWg4o
xpeGkCLqM7qHFBjVVhPt1AfmdklzmVx+p1KH8FpZIxpB59zjWvrZ9JbwRvp1jB/DV+4tOyQqmscI
wQ34SoEhAGeZ4zNVIGbVwaIMTGyXxR9LkIgvTk5AYFEDug3Y6JJCu7RryyIXia0mJtI7nOSiFCk+
RYTyrFPZ8JAydC56z7oFKhL6TH61sfH/Tq+/LGviY47zEx57Gq6tbJaQfQjlP5NB6QxxaBFgcE7r
bMdscmBhePiLnWuCMtnYZcH9ozrphy2CGZOmksJTtKF0PDyO1BhQp6UT9KLjlpi+5VWvaGwBMMYv
hYdIFBq+HsSjW49UyA9fO8nUzBTxuRrZtcvE5SzNDvvVSsXpEWE4q3isabUatvI6Jt3T9XNdr32i
BKCIOch0N/WojxqPIamNQlo2kD5gkXCens/HCxNzo1wJU/3TzMq0DkXW7QXzBCIipxt4IEgFJeTz
9e3I9ZQaelJS02PO6ZnfdYjKDQXuAAVgct8m2FaFedsUiz2IDHQgOngERCfwy366mpk5kWoouwuH
AEKe3MZ7XwtZU1cEPT3EFiIEIx19xvhj1k9jMolZWfzHNA85VLoaD8VspzpE4Hk4DwzkxgMqmIuJ
vSCAcULfhfz7INvWIi67iQmG27tJaX37uBkhKLLo/leLc0qLOfiX3EtlM4jYkye0HlpYK/06bQoo
1dn+gL1tw98ktW/QVzr7lxfzFwB7TeMha9Pm/mYCysLtjKnh6Th9+G4PvJuADJJOoiGdHjRMY2Px
e9gmJ+7Xa+5cnh14hxC9aauyc4i9DZNz12Ku5vhVnvs8wpjZYx+cN0QVRBQVFIzsJINEgOySd7sj
8W6as2sihouHJja0CbYUwnF3v7eRG46ar7Pda5blyEk2bN+CRimSpvznBCMICgEya5BMufPT0A/F
gwKPQdLmdbv+DBT0oW8/PY+67aNlvoZR10JLj/9DUfo8+FzOXq0r1zP31/w2U1PbHfPtD9rRy+Ad
Bt0N+KqBwydApfCOc6R7CU2bQa8VkTRUVani7aBuiU4qzWm4ypFOpO9lXcMwOiPNRS8FDlRyyj64
p3mSCT9CmJWMH5wfcLlkLW7KeyYElvpJZfR99maSmHClf9L14ztKbw1sf7YCQcOOsSxK/lfiB9Dw
rcBso/DnNK8Am7eccWrFRXnsyLIclUzkMhggPRCJ1QSb1x6dP94fT3GspHbvQZSb6S4q1Y/gt4+F
nikrKc8pU8KpD3LsKKaLPd7l9I/aeExJ5LmMQNhXy6LPgwIhHufQYkK0MsJOYxn5vEITZCI+x2rE
LH7VMyNM9lh91pmPoAeNbks2GZ9c1I5qiVn77ae6hsUoFRmYN2x9tHNuxF5TLKOZLPLvPBZSwl2J
TqqQXg8ke8AXbKQipEP7Mil6Vqr+YMFzn4AVQeOPwaNatvIEC4lUavUcJCEnELPD/8nhXyX/Mrpa
SIohZ9mWCFW896aaKqC5Z4alaM9lYss9dGAf/QXYgVviLusmbR7MxSXZp84XN0yyuXejyQvNQ7OD
KDYtIMZ4EeAnHdBOfZJ/brQshSPUMMRe66h6bJJw4yYxYHBB87Uz3TbeGjirVJQKHMJqcGv4gZJR
8zct5qHGeF8rtLoZTlQk+CtYAagAi3OClhfTv6e9s2BboBKx039anaRZ6kf4sCdfb+FW2X0roFl6
lp2kbXk9YERERXMpqgxG0KHIq8+FOIpRewA+tbUwoCh7V8VqS5A4WSGeULE7M+LYyZTURdNB8oPj
f+JkkWG0YCk8Y7AA4noH8PwDJwhIIsXpH3cik8ERZ35WJDCn+UauixiJKm6gIXbZAvpuipTFz1mS
eOTMDUnqlblux8KMbgSEhZz/iVTn1Fu/SROeld8YGBQhWsIRHok9SUNbCCqp9QKJcEwtG+BLdgaf
DAiQzlqULGpWIjrsdMroDxCXKg1i7xfIZdVoPS4QdSGf6V4WFFSkh6bAku4Gz26VU3JXqWK4p0ny
gmgSQhbYe9a1XGX12D/9zYFwosh7Y/fp4SqEeIQZaLTUBVTuOWtyJFec9PME3Y7eWwy0rulbBFHn
qoqKdzjAi47WqCZauew0d1Rm38se6bYwxyy4pYUrrLCXbeLe3KAJX+60Af8Uh3wBLp/FqmclQKIt
nZfA6lKGODX/e6zpCepEzx0hR6FrmYo3RDTsAZXn5b3FDTrX9D/AViU/rd48dS3vml4edxWx84K3
3FHRdZe5fSyveYt3T1dSPRSVMJ9NSDfyVfkTaL0paGPnb0kk280MY5oJy3yAqk10qNWxaIDh3awu
rH5GzjUeKDOXnuwxb5U0WPq4GNCWxxD3SQiXUXY8WRu2XKTS9kYiXJNE5hKZYvzTMmioWw1KmYUv
6Q9tkgBrNZEHqZBXeHBz37YfDG5nUwtfmykqcolog8HumTUd437AFg/QmObBFLweK+AxgWmyGMPj
tbTy/DHhM7q4JHV6uIUTSyJIeJHm/1jeDwzEYaXXZFPqeTX0erH47/EmdJGRV/uk7xDMJ253wnYR
DTtRJVDv8IKpN6ND/Wm/bE1HOSBcZUGPvIbz0bavT5/szBMEycOB5UP44l2+q+PvPXzxKNIEt3eN
11gwgmgGo+WQGidqxiGPf5D2LzUxUQCVZ02mC+ImpqRAgzIAb30p4UVgS6Yt5H0bw/EDzhv41uiC
piikzlcVAjNTDuGnhQq1dGOZwN5rC+Jddqchkf9vq48i9FQKsEFcsbJIwXXUeq5Bnc7iXMW8ZEph
a2QKgbLjag9GFCLt08CLevaBUt0sW0zfjFwuJlfKihOAqwYFR9Vb5QPZdq5psFnG+iVyUCz7Vqh5
MGKislVQctBCUq1htGbxVpj+VfzaBsUUllSd68qFPCPM6E/2lrbFbtRrxLKvwtyL30ySn9k+4Lir
nomeaNugDE2B8TM/mlabLi4Ur+nPCRm4lkJHUDRYUG6s0ZEauoXl/CqS7b9v0023QHSK3RTGv1Zc
G1LAeSDr/YgKoph37FYxpqBIgJ2Md5eKH+eldBv+gjdFbnx5vbWelxic2ab87132pGRN+Few7vZ4
+I9+FmYK6VAM5S+5ZYWs7BtIY9iZ4WObfq8fQdhniQAaduBwPXdIlsmX7eUYwKFi7Uf/Gap9Z1Dt
Bw2rznyH+aSg6HiHIhFBtnn1WScLQ7qSVrzuKq44HyUwl+3sV7JU0P7mRNWwY2PH5RSmOD3zMsad
8aYwfYDDgEKwq+1/T1oAd0Mb+8ZDhPHlmyAPaQP20o813uamtkKD2I2njw+uX/hCEqBDrrt6HBA8
P/vl4roqs81LsDal6fumsc1w8XdxwVxEs3b8XENiBmEiK7oMRV1tdXsLRnaiWbHVy/EonpZRORC2
ixK1joWfLdyJx30FmXumSiQZFCrfXFKrLrYMyA6nvZLXzpXfQKxeyDNeNsKR4POKpPkVqQRZ2t8L
/RuKBJKoXuy7Q+b5wCxAF7tw4yMQD1PmdLD+wfx8EiHMAYub8Ou7BJF95lyxWHFb5eBU6WokQChG
Vu5/YWszN5zKJM+gOugTjrJxmhEzOmA8cN21nvVW2aDZEjdtOyHeJrhtV8Q2VAM3J5rMbDnG5YXf
uKvlYTTQRHWU0Ti9K98EbyiNRb2nrA6Lq4eLa5i7esp4eKA3E1xUC+ePAzHbPUHYnuuIuErPtTov
CB+nbQlmhr/CboWIjVRYcnCsNoANXzwU7nnw34k1nz4h5cwH5AogdPzQ/2bu1O95Wa31KTdySEbH
T8UscDFtbce48cnZmLrBkAnZNWkvQi2GQQPXUzWqAu2H/p61jrxJD2jPG6svAh/C9koPOXXeeK95
41hRCCdI2jat3kjddceZy1/tJwKYTTSm0tLQmZGV6lR7EdRnwAJo/hhcE/OUVL5raJVsrEWXGb2M
qHEHcx4fJ6mNIOmVfbBXFSn9q8zEfklDL/1xW6Aw2gSwUazEED0CA5j/2JnNyQrqIJ/oMbvwyAN5
zTgbWumx+fIOfEk/iBmP6xET0tY+V6PMI/S+aDFDyKi2YNb/NFY93PyhLtMzDqXetAxxgCSjclUP
CtGJQvuBGGI31Dh/pmMdQd6h+DL+LgOUBWV9TUIlORfldXesseiH53uPOoBVoieJYOILjc8shrcK
kfx0w2j8Y4fyPgoGDytDRR7D8jHCKr9xM+Xybd47kBI7vk1nHeIknN+sNhd40uBR2YITB9YvZHp6
46kSstzmHWfyCyGZ2VtchPKlvKOLr23paPj4mWoOQ/DGM8xzYJwFENTjevVRa685DHIpjoO3wJJo
dq/Vlq79mmFhl7yL/qWWnep5r79sDGzumuTbC5L4u6QxW5VzI2vEsJy5VHZeNe4jtNJFgOJkLwKm
vht9oEyQQPordFDVT8Cj2tl/eUafe/W7jHCvo0UaZfeCXgZjnJAuF4n1jtfmfZhZP89BxYt6m7Ml
TOEMXCG7jnfk+Nhiza1E/UywS0KvUgto0xuGZ+TKtoiO1Lsgi31mvyfI4lNNa2C0t2LKW3z3EVAp
kv6+cFuz+0NDGJQ3I2s9HSOhFX+QR1TTUHj9pxUJ0ypVuu06M1BrfPprD9ebG0KDKpDFT8J4yuJW
miMr5F+qSKmlcMcXwaNk6sdQ1omKe32+3nvocAP3WvfbPIDJF4abiaNrQa41GxjBlvpyBKFA6Igi
vtEl2uFLpQ48FsgDtxnL/uHjbtXC6IGorbql9Ynji44T1Wzo41w6J41tVzCld/OYxRprhHPW8fzF
DRhh1tNJT3gSz+Alvfy9I3P6ztR4BgN9ahX2oaA2od7q6pCmwmus6SmDSVx8SZg4tL7vYoatTzgJ
GZdazBLermCqwXhWJzA9x+nx3X+4ch+XuyIg3qaol6CYl+p8KnsowffuSfWfrAhceowYNnAf1Oi4
8utTH5MINwKHSMMBRTML0u7o3JJuiPdGlmJPpf8lwLSrkIKAZ3WjEEU/TuCAzwPtSWJeBDrT13mx
uw6NzLEoruzZR01542QFv+jIqNExeyu0MvAc/BVWw16qS8xKZmgpdjbAIaHCKVwdm53vOclMJgUj
FrJFaoPOSlWX9dtsemkuX7VEgMOoudp5WAXwdoXA9MFGwDXXx3PzZtKSfXQQrxoR1XFq/s+I07vl
N18KuxePK4tRmGu/ReYv7UqXJ4heFEq4uoFCRw3EUAyefOy27xjBjYS7B0I/Ac5PIuEtKM6CcdW5
IL69lVr/VO6q+WIVzyweJQM6lA4vOTXPV81UOzi6ejSP3stuffZ1VTbFgtOVBjTNYhn4wwy0bf42
S+00sNNavkLDhIXsNMHlIZHLFMz49MNZaapFccBnH9o+tVryytL6H07CY30nhuYR57pX7rg38QQm
QCy2ntcOVS7eDH+M9uNVUqQzEcO3chnPmKmOHv8NzA/xXK3AR6j1JEav8W0QCmOKz+bIdtGqGu9U
jLijRf3hEZ7AjFop3unOKFLe/Zkk2L2smFWRwADWT174C9XbHyRtpIs1mCk1YbQwtrlP4JKBKjxt
7O/PR+lWQNTBleiot3kXT7FzIzSRLMoSAw7mrGU9Mcf5+TzSrhTCOOTZfmh7vWwRbR3kSGRSJXFf
EDWn2ZK8HFMTMkacW88nWZ0vTf8KX8wfYqDCCAVrILLPEvuP3XgcT2ezXwhur+hQq84u9Yu/8cl1
Fw05Rg71/23//WECbqhXuXJr1XfLgRWo0woh9JUrItnk7b31fr5O09CD+iH3CvfXc3AR/RQUWApQ
ybiS/dyJIH+0Xr8ftAESHHOAbg85bfWYVCxUd/MRbRfpnhLXcEL3TQY/ARxoO37tlP0InC0T2jqL
fAkCu424XgE+GYbcowtvAuwzynUUbN5FL4ZDTmVdiWITKKrdDNv5A/yqkj/bt3ZnVgbIcY87ixsC
3ooduhQuiNcQvqZ3VmNFPajY+KlqBXklyUOA5Zf37HX8rHieQ9h0KtW/ZFEafOopbg2ELmS603+j
y8DDE+rGFo3zn2j/9QeV5+9zJNl+xsHEtWegcOHGcziSsSZsrbBUkcjhits1m1v4CF6K8nFgvQOx
BPN4d2R6CsY8G7KKw9ISXYsdR1b2qIPKCpATTn/k6KYag05g3NXU6ysHrAXoiW4Wy1dZyZ5CrUGm
tTc9CI6VPTscwspQt/qE+YZOAGzTnxRb84o87A8dL0DsaH/ILqyGCKGloX1gtUIsvB1GArY5AAuF
EDq3KzRYr/pbz2ssRExOxAGj3A0DDX5cY6zE+NzJdEczZkZdO/g08mo+eDvprxPwQUg3gSMKKOhz
TEB8UCLAy78Iu4+KzVjPoQNC7dTdUWsIb4D+OjydzJpuSyM8RE+VA8Lepb4NUMIIE34/GrsExz8Q
M+AeD4cVxpU3YYuF6hr5PwFJPDJxWXWDIOogM6bEz+jSBMmhLAimWcZ0eKcuIZNnr8Hq6RD4x1oF
IUU0Qzrl2YDaLvsCPWtDaKA1GWbrFbYVusWxO50FRlubTG460eDNuE75H+/iA59CtDsn+qUAAvmy
daxEDxwiij/w9CqLol5o6uqoZ34QqCCI9LRPxOTOM8N27LvYV3FvUaNoi+lhF/ht7PlP9eYV6CpM
jDQ+WYfs/w6i3talCLyjiltLTfM+E3a9WeuNkXijTduDK0Mv2uYaeoylr8Lv7RvH2nGvjB/8eWQE
S3CU5/KNqVZAPG/lUnm9RWb5DCRte27FHB+VgxQS2seb9m7wJuRk1bnnt9hVk2onbFP4M+kNjUat
F4019jUwC1w3XN3RxeHnmZcj+AR26UVgkTZuiABBm2lYRbEX6BT54qDT0BSC8il25Ipfdk9WJQjP
04RKAXI0DGXCDpWZCnlGZeHpTSxVlXcfrZdK4GZNRQrmTyG773fEjWYQAToY3gaP9uaLP2nWSEwR
LfQp/I4HHyBXl0+7eWAIYtq7f4/PCW3G3ZkxrKKQ2uN04oRbBTuEc8ckIFoa20E68B7IashhAczs
/ct+Ft9xenA8jtnJPYn0k47D0EzFwr2M0hxctJoyuhuhPOsn9Xk9+Zd/uAGuXGXhBeesj8WiDyeb
zifojADN+z4qrDvtrG56hCQmKgL+jYazMymahWr2fh+Qvf795QM2rDyJjavrqbyeCnOZqNzU2anI
prKbwtwpyyaitbdToISIy+u0IAb3XdteiOqxE0JNgwH36lC/Jm/wZ1Irqr221LaBrLyJMDhNJghl
j62Ch1wflwho/1iyGPbhQM4Xj00WAtrcLUTNRI6W4w/L2pGQu5atd2JmV1DUgaNSSply0mJPnAzE
yy6sVztAkHttvYR3MkKX3NMLNtDBSZWLjKis9pE9gQ9ANBWZ9dv0xudTppFQfXIvXgkqvyDCyPui
4LOa9+NlR3hPluiSIcS/4TOlM+5n98P+ix7bXph6HYjdy8xHWivUugn3MU4+GV2agO+Lj03zQsLr
MRv8NNPvGkJv3gx+9mrEBwyFSLVwB7oZSBQGkImCc4pDlaS0o9/h7oCjOEqrjSDUVLvpQ2aWZ+E8
2kUfw/c/OztAGE1EL46GBcjh5A4d4I2SrAaqmXV9Svwf+WD46Kh7DoQvKv5tFBl9QZmPFXAT5KWx
ga8oUmL9u7SDUUoXtEphzpSXJERD1p5lVCHt5VzuEh5MYfWMzUKr0+YXjYidp2yZjptslJ7+TWdq
5OKw1xvbFIya2oFYNtck6SbhXo0Nht+rP0+yv8sptSK3MbUY3laiEkZTZtjl6O9OZ/0pPVh8jtpT
3fSWlP4xdEbP9I7ydfhKW4t3sCJypEgOIsrDiOR/dPfLS3svW+mAfnc2LYWe0/8NGzi0UM1d8nhG
Yy2ZkvfuJU+46x/9dS8roRlHBTwjX3yAdL1ISC6DegqMG8/gcDHj3SccDJQ0VjZmzin+R3r7F05J
wzLy1svafDJvmcBj6uh5DGeVI5W6c5CX+I4wtHx6t63G0NX9TqmNIx8sj5TMTX4fahDy1RJldauH
gykk2YErqb9za1kYal+Wau6ih+nw10p5GbTBKLTjVTwoP2X79KC0+6pqcG7aJKQiw4PzjtzrXJsC
BHIqysDBjeh3OoMGsJgIhrmlxexN1O0kNDzsqUzpIAVEGfICi9AMXeNmVCoS4Qn7IDHmS81dTrRB
E39ZbrLK7mQBAUhh/Qig2kxulCtPZ58XmyfyCW/LZe2/6ZwHAQELcEPfYfS8Yh18XkP0aqTouhs7
6UQWlW+VMzvL9FQKdqaVnAPda+FtOZLeZvZyJLQ6kqlDNlOUiCfGUVAZ/NwrudESq9NFpvU2Othl
kM7Hg9/DEdwvqplU3AQuWSHuFNclwvio08zfOkxkmB7OoVNJhAiSJVfNJBVAMpEFzkQ5cuosjCWY
9Bx7/SfFz74R4AHMlH3nCKO3kC/xLzzoS46cKs9ZR34Qq7enmAi3ju6sycebcdYBdazveoFVpllm
KqbHu/QjgyEw7YX1Mk6+QAF7wHprCJgX04SF96K9z1eCvnXgQAbYiIjalcTEd0MOOIcHWXoVULTe
TdraNe9L4UjVTNBvMRKAcUfSXDkEcXxcY5lIATkSXhGpnUp7Wv8xi4Srb+ypsX31OBFDWt9WePpy
qwZ5xINopWL6zJ+e7Iz3GJOZTeWQenBHwziwVnyYuymuSOu2adIjtpEBMImgDfxt1v9IRse8Fs/O
yHygaq7dsvUg8vdA3H18YAntptILCfS0pM1RKilidRdGohVnGNbCbV58kqPex2O31MGvfrUAmZ1a
l8VP6Rwitq20pJQTDh/niYylC1SguEymjgqv/uox4Cp3mcai5unPf35OoZCNMRh60s1eB07pvBYK
nOqL4k8FfQWb6jvx5h2zA3UsgEKG7hOsNhTfP5/bqcUnanf3Hm0Dh6A/7BBiD6Q6nt7bntE2TwiQ
lAMqJdDkPQJo2jwm3SK4tVfUNbRKH80WRrBKhKze3Xs49omtlGK7J0JEzRmUEC+jLfF/RIW56FdS
mW5oWbnKGt+iz9mZy6RzS5poazxjX5MnZ7WX1KUPSUWKbZHbPfD65adEXpmo6NG5LpsRmf7SHhye
wjdZrPPSTnrDAPeV6FiC7aOIQzswC2wPjifVJquyd0ld+qTPRmQfxJX5fn7E/45fV63OMU72UkNM
MFGanlbpA8KW95Y1YMOYkugXiFiTG1Ez36wL6MEoQQPEL2MoaThER3SFDdTEVRebUEDf1TCCEgSW
Qs9pa4kk+oOAkTnCtc/VHRx38nGTqmLXTpGGOo5s0Wh6p7SGLlv16dtDjOPmWWWhlFw0NZBfaTAc
3ihCSidhkhFZdvp+NXvHZswqeNHG44+Ly6E3ZiymQsh5d0RShoa8IvxmTtrRHc8/8Xzuk77/1EMu
GL6GvKAM35P6dyzaA3oAtGOOK0EHvEH9ErZMgyj1FaBYXtjBevbh9V8QBAXzxNQJ2Ff+3694oM5L
z17fyf5ABBr42+gukmiLRJXbaYx2R/zvMUYHUYQtPcVDKtB/p+db55lrOSktdoUwhKNlFYX/6BL7
wDLeyCCQ7BG7rgDjveA9eu7n1Za3rfnpcVj/JE4w0HxFstTGKQIkSx9daiNFQitpHvRD32e03KN/
H+XLyaE5rYKBebVYneWJA36CLOXIdlW65TPvZdptCXQ7cGwJKwP6104gnL5XAck+iIA58tXZ1csf
Qqz2Sz1GA5Wm/0224MvnapSQfmFeEqB7+QB8oVlaKKzQo4LBiLmG/7X3kqUrOuvTYyYgv4fPDnNR
rDNdVQtqfl/MfEN001yzP1D8Du0qjz7sKI4FwTWXuN8fjcm2M1+bud9Fxa1qq8HA9hhPJtHTGBpn
52LkKpCIV/GaAIcUm8ndKwcukA7Ha6M3gFIJPVWOgJqPycTsvxj48rxo26ieyqLK2+fkzXFwYZ1X
tf8l8RrbgVWjZjNg6IsL0KxsMaplJtihbvMojAnkBayCx9hLVHyqhZajWeo5mvToI6mogjl1UmQK
+2linNlVtTSSAKHbAxFKGZj5b8NGCeUProOuiKZ/sg9gGu/a82hkJCofdVOOWzk16GpyXpUIhI6B
lOckkJEfY9eX5Ale0UvUTGbhXHHMGunP9AmwcI+lQUMCdS56uoU3/lnuhgGBQir75ENgo/IcI+q8
gEsu/210gPi+54t2g6FvFHNz5dR+0CsicZ6I8lOl5DYiyDZsf5jkMo1vQc1kyvEMFifK8IpCyonM
4E0tcP6TgJC5mqGrmEHIGpLSfm6h2ZrSJFZq9/2zT7C2ynJO9NreZEWzv3q3o2FuNM58afbUMWqq
sebrUhh0Y1lXW2MrxYEwtlHRZ+hz5Es9hAAiBJ8NvTCYXLY0MmNxYdcB925hy+tOelG0zn74h0cX
sDtMO3KQTt5xR60w5Qjo+9DczqxjBGpDcP80YDR13EqL+jGeNnCwisgZkKWsrfrvaPIKLbRHjoJD
Y6po+xAenR9WwLbfElVU8h8PoBWS+g+h8Dm0TzhkcdWRTlllaNZ/77HUZXnuGwAdc42EllbiHirR
DDjV9uP1yOlNKA1OMeYppbz6wm9GVgakrBuww8BvxUR+aPOArynPmVPTf3Kijac7UVz7RsQxSaQO
UkBhZZYqeseff5XRbhA/PO0kfY6FnGDLijNwuzduKiGT9PAV6yIikI6S0KjaeJE31Fcfgm0LANLQ
yYJAMNDRSU7FwCQ5lkOYdrS8WztAfxDbIiVG6lA9YyY8rA73lEtFPDOcPeWoiDEF6xSUHUvGvdKG
Hl588dbViL2l5HW+lcurb06yF2nVJyiP9axbuqvOzXvJqZGpzac56d1YcKEviuDecENuElo57wBI
zRhl5V0LjHHiMbQB9LyCzGLTbNSAU6xlvDUzodWFPYHdM2nXhsrnKsH0Tgfy+y3ijZkYx3pcnS0b
72CpNzRMMFqC6nGdVGC+V7bOU5jaCMinbsNT+yepvENBZW7JZG/szHasu+9Ag/LLkEzpcXUhQ8Ev
80EOlOqrLVcXe9XMRql6LkXflE2LtGia0fG9mc4HOvnAOPFPzoXDELlT9Ld5nJFzmRdp8Sl2xx1l
kmDbSCa3Up1RrWlp1mDSD8cYKv3FhlAXIAcgzy7j8K2qoqTxsWdHHYjLcJDLyv0bfpG1G62KA1HO
pA6ITLNb2QkZlKNVjekwIgW/0ntHJ4CPBO6ty27Pdqd2429cTQsUPcyrUzielkPpFy1OD7Spf7zd
W37iIBmlVc+uGQnvR2bG9zHq1JyVM6hQ6oJnLndAZqXzcYoUNjI/q/HUn+6EeNbAtIflPEliQH/c
uKcsWnSy+FFFzh0WEiIQG9MDs57v38xHTqeIULcdth2jSpmpyXpa6Oc/pbyJLY7Mbbem542GUDgM
XdyaW3YnEkbnXPXY1womxq54U+8a6954f7Hc98yKJ/tzbkXIc3MO5x3faFO9rh57QvQA569iZV2K
/ajZySmewPIOFRnAhzhNTVq80C3HzrqsG/A8kH7eXTvC50Id1h+zUtb7Ggh1GVIjfckJoBYWROku
rVn9QsL+KJT1zDurwdxvXvvtWFIngztdRC3oqxlXFtDg5Ou/4qsVy/m+JogkOgd4wZ88hQqD5k3d
+WdAJb04UJXsV2RNKVx/rbtcrT29ldgPhxKr9/BuWwtaTt3GfCcQSO6QRpMfu0s3TUdAvbXSpRlQ
qsbhjT3Y5k6wN5Ea8IgZFKRNN0U0e1erQRzemO36cIJeIcrDSDtJTewUmoeU5QE7wkhVkrWaBe9K
IQ7zqPBQA6Gwe9a9XLfIVGw82IyYbLT2ebTPlmr8QRf81kbAq7vgiDNlUNSg8srfkmp653qe8Wud
I3zQm+6rrIxXsJkYtN/f/0PwD4T8hcMxlQHfGJVA4hshMf5ErraecRs/GGv/dzHdvcIBENHT8J0D
BDvXVabwq2WWxNOf8xpfxBsMipNMX6++im4zQrb4SFCLjtdaDueWr4kH20sK8RtMeu1sPWJyzpde
5QsO1iCiB+iJkDsZGX27NPLPxfoaMTr4eGecn8c8/7Lw8z5L/4q/1jzmN4eh0K4N7xvoX/0xDA2b
B8U3J4x09kkWvAHSTQGPQMwdLpwHlS998p1VIcgb47JbK2B80cdeIRDNGlE/Qy1h8+1eoa/OlSm8
11UG+xEM83+7iIR7p1MGBgSXOhxOj70wFnpCle3Q8aC8My/bVIWyPauY8314BxAwNTfOILr6gBSE
c0cXxfW+1QPmzeLDUiK3M7nA4zPQ9DwQNy8bEKStMZxzgrccQacxtzAqJbxum4XfXKhGfiZqyY2X
wZpb/4gQj13h4Zc7awKGRV5TSy03nB/vS69/CkUsAF4dzq9Ycsu0TYT2AS0SqDSRzzGchoUX9Sy6
QWKCnYpOFK+nyQAiSFjuAC2Rc3zbAVaplcmlK3oi8+XHKhsGClncu09TK3NNkViyAKSh7YhuX6Jh
4RS1lX6qIfsV1Cf9ddlhjmPbIahWFh8AMEqIhT7Wg0y8W4ZXEeHKVLGJeCmctWh46ZE5MuojeA42
QBcosdr7gUoY10aLwDQv+CkxZLudVNFziftpjMRB66HRBeVmkiOecdgfO0QbeGnOuQEA5Nf5JlJl
jIuOiJRM1ANn/fTaj3tQEfFGanYWtIUymb1K2Pz2Wvf/wTnVNr0H33L75y4noWo/PWpC13cmf+wv
HilsuzB+VNPhpgPEXQQ+bfHW/PhnbbuYhFwokytAjVR79eZ/TCBBWUE0gVySQfG0xI/rEg2RVf1+
YM1mW4RrgSxuirwd/iCd+Gudpue187OhxOIOGRrPP3hIBURNbma9p8tLsj5cDJJGduufb/wOVnkH
y3m6q4n8DYGrMEdNpugvC3cLEp5oxhzUIxkU9e0KSw2gE7rZ89Lfy8shwZ58mXadskEBCneLyAbQ
4kKeQBZbYmIesQ4YTqH0BuXTapoCkJ8zp0L/skEuwwUvjz5APXWKjDnnL7x+wq18EtrW/O8thsLa
irEpyB09ZT6viiolOq8YaQ/ticd1qJW5+swYkZM0A1hAFXF8ba3qKf6P8rxjtxwWMETzJdz88HlX
NpdNXQkX6oH4Rcz8LczJr0HQtF1hxow1FewzBubexobKMiAURMoqNQYx7RFM/nQgdw/P4/iEqsue
CpbrLqsVoROxzNL67sjLi4MXMniIxIBuEpPQDdM+iLTsXRqeXKvEjC329e4x8N0x0alK2WkQ9CZy
rpqaqxbibloG6FirVzgsM8V3nadUIEQiliuPm9s65pQonCO2h6ZaoK8Oe1HBbGx20PD+oUV2hyJw
N+JGqBZBY9VAY5EAsahyChcy11GEC7LTF0YX6J4WcYA2ojBFS3l4C3jdI86i30kgqdK+CkYiZP7e
dDcxCxECzhkFn5jGNU/o6XuBuV0HBkdO+ue2C1JQ2z0wutIlBW/iT0h6W5CoxxLRzJGclTuwBphy
yJIHjDg4G0Dd+vbBZJDvY3nWYLQ+SHRLy/UDUlzfyuo7PP8DaJRmbKNwYr8qOESVy0OTPT1XOAA2
smbNPaaluuSglJaHUfXPMeg93+HodkRnjvfUPi+r5Ko/2KpiEnJW4pLSYmsRpN8UULiGSzTH6wvB
uQhM+CuoGYZvL72d5/zcCZgzOpF9KVdv7Q+Ws8VoFAPic5VTio2X0+XSEvAVo9snmCk9RDM5Bs53
qeWjCV6osmcKmP4pNm4yDLXLy+AbOk/3V4w02MOKLJ8ibSX58fsnNMWsslS9I2PPgSbr0tI5mO3b
DDnXfJFDel/g50GGyLB6AMhXnviAxZ82+lCJtpI1M7QeWhpegPHUGZjJ8EWpwnIBldNsp/JNyykW
Ch9sWUKAUxLe942bppL5oUR6suhO8h4x3vFB9p4ueVcVlAdFmeM0Fl3PGbACV7f3k5KssjMoUxls
Eh3YeRO4+bW8cFiwVi/tZW76XAezz8MO/fStUjUtI0Gdq0IAOql2qdfTVGuNBqeFmJ3UODSsNulO
WQo3BXVM7pLVN4YscmzTyCVQMXPRVpbut/rOsm7dBrYOYLlbdf9MN3ZphtpNhIyzzSVgMhmWH/K9
mPDgdQJAPafFEZCDNnTVEI8G07kZB1Rn742mZgWVjO5xXYR/I/TjsghAL+LbDj+6g5P+/213i4Yt
KmiY23q67+dM0cXUN4Pm39tq0DjZxCqfYCI5t1d2CtCTWQ74aP+n3rTxNs1BQZz0ZBBit3uldJVE
cI/vkMt6FOyJhJZUp06rnExrlmoeX0YMIeCaroaTaxnPjl0/0+yT6jafJbMOTil59n0oBcjVI9I0
kYLu06FqRVL3UT4rbMp1ig1HHp5PLo9hA7F70AwltXc3lkNCvdpfHVKHLrY3hoV0SQ2wGVwogC0b
AKL7WYvlKlA00jiUOaN1P/poPLincEMlNjckbORksQQXbBEcd1EVTGLUmGf9BFzctRbLu6++0lc1
P16GNyk2tmR0zaENIoZJXkX3zVWwuGp3Wqd2LJDBWECSWquzIU1FUr5yPqTtBZw7Pjmw/Mr2CjcP
ytV8HYkBKJ6Hq9iZD0mUUZ8JO7lIQZHD6UvcjW3YIhNjA9232LThyPrCzbj4yAymQFZGluerSE67
5IzfYN1mlHDYN7LeCu9D1Z8W3aVrw+t9tuz+kgj0vcooAqOqgpmpMrPKGAg7OYwo3MzWZQVLJlbt
NEWF3MR+sT/1MRvHRcZRCFJQaOAyyAsSW1hCmQBr5hVoXrLWbEhcKCDOjn29P2WZHV6jhfrbfEOj
NS0+8ewq3t80yOt5ysZhchxiGCOdmW2O4t2IkXWbIbfhXu+SoTlNuo29cvIEh4nuUFBSUMvSKWmD
MIRZzZB+YTgi1q9xInbnfvUgiv9VMMKHxXmvuW0n6+5/q6r2gGCJNVy7uENgjdbBZ74gTkISubxZ
hBuLUAPZ/UBZbYbn6sYAk95eIo+y/240hxWHfFVfJxvkSIjvMW6dSlJpFZ2+BScVguU88PjbeXy7
U04QG/YmeCW3jaJMTOsCRbNiqfPmoedWMfdQHg9cNdW6A8+ibFkCmM27c6DsZckGtVDd9pbnJVt3
sKUPfmiR0XTWw1+MVEN9ngvU4Fsv9V+Xh9n6gx+v1jw1EOe6Oc3Zi4hd1zR0x/MsHKYCgWIEdwbz
suWLLGhGTSJ4RmDzjBITZXWsEwLsE5SLJ/KXG5dSiwNKqGnHdJL1bF615Vt3Z3UbPm3DJ2CqOmEl
ycY5DhQ3CumUZRzXROdRLjzTtqZoyprBvCqIQBG+z3s6s549ea6GwzG2dYcYy+4o/0+DGzyUWbOB
F86jiQhhDbXtKpOqgrpBJCLJqqY2h8z8cZWrfVforBZQ80fY3aJbX03JCTfi9qb6X8hRi+KVJZ1h
omyZycRHw6YSmY2Im34yQPg+YUBoLRiw39S3pUHWOhnQKUKYjWfwVlX2G3jZ64mqf2iRKbMvDG8i
J1q5qyUBarOPfg51JuRO01sTJtCUmnpsicDHKU4Sorxr0+c0UYHjX/ELk5L9i2S1R+Z1D8LsJNSl
vBnO4jpDWROMEnc39Lq6B9Kbx6sPqrEb4o51zldKBbiTUXd4v2AQPJX7NpxKJ+djXMtpduG///wE
2PL5BM5nog5FYQGFZcgmwD1iMEErPYeJnRarr8QI5bFu8LehYHE/foyl7fYytBCEBTwGjEUJC62a
CpYGknvFrrHRZUlqy50Dd2IxVY/Dc0wSGBEgs1IE9W9U/dF1aUEWN9DmvaMl4QKj3fKMVbArlW1L
ddX/krhXceR70Cu0Oy6OwluU3uFbW3jMbjrigoYMCZ+movOOHguJJf0XyqsBKYPTVURtFVr1qtqa
/Giaucfio39mnDVXmnvUOiCIeW26LGJsxrVoWo4HGNCsK6YhmZxtGwWnB4tAp4MyjdnEOFKCcH1S
rIQg0hnNcJXQjroKEZ7t+LYBSUrbrKX3/P5oGSqVdR5N0+Hu2A6uFOCIJaV/3YXjfovZADvuBsFT
5XNDI+isPnSA9f6XQBjQDBjmioeAjPRZdvHb30obYNxVZcxXN+5QFndJqgHUIS2kP5Nr+D8tbGjE
k5mDZqG1F7g5dNThmABveVyx14KtVwNLL6pyNbbyy4m52uxZBLBgrhTtNXTrx0O7HAvpCr34eAng
UWKdv+7CTm7khAwpEjl67wI8Tlaku/UKAh72IipHJukU4Rga8g7Z206MgVbhImZ66G4cOHKljtw0
Rru6LG2b2covCwNm9d+0GxLACOX4iaWC9TElstRWnr021+21JtyTYNG1awa9ioMlF2OWlV5Gmz47
csqxw0oqaOiAlpnQNA4ZFcwkwUrWQf9wTvYv/YOjGRNmNySJIBmwPFxx0v+UItIC8BSqzoJ4c/x8
AG4rUxJ4EalrHDGwt+cqJo1TQ/IrC7SiPsGb8TC6J9wJQdsww0vS2reEMcb/p1GPSvjUwgIVTKcO
jm6zN/lVFiPnr+UjSDtZGrlHU3YttaeLIqnkc+YNbPPB5aPDp7anxOa4+cviMwSeOqiwvA3MhheF
Whg620lkk8zLHKZpgVsfC7lxOGyc1a5EOgDMK5LRboumpMkzg1l9RG3xeGsNr3X5Di2E6bE2fGSV
Ga8w/hjAmpuRfQNm3pgGCF3LSfqF7zOnxUfgqT51+avDqvMNgXgyXFYvNvaKCQIKrNrQLzEpfK7D
sqqPObnYIQXCx1DIg1X2dkhzZIxCjl2+Hj3WNoh5e0bkH3UDLq9vMEVBRe04oQgmtpzcZM6nFfEc
c3ss9k0hmO/pN8egxWJ1g7CmcjsYNbmijEiSfvsOb1Mv3JbtaRDAm2dTXuC941/PK30U/T8N8N6O
dsdpZKwP5LYhnYwTNTk2G5qms492dZk6qCTWJ/Qiq3gwDdNVZ1Rvy67cVGhhhAouQCyAJYGcAs3X
5r/WQUFWjrGLI1j63XpivX2CXduuS3lJ1wHJI1jjtJ/HYIx4g/qVjvHG4D0xxrBdMqa2y49n3svD
cBzHjwdBReBM29Cs3CYkBzKAGybWnTs5S3kdNuJKn1r6tNKBiDgM7DFwKBj8WUoLe9vof/6dtRfY
/RTbcaET9+h4AOXmA18SZ4X9pqFdhmSedFalhpwbWMriDGGXdgKeAmu5YhqBFBAhqKwiOJcW7q8S
7C5KD6ybLCNqY8HBHcFyi71rko78rhXJmsytFFw3DFoUyTjRpEGMooJfczizfO7iCm4yFPgXxwQR
AKqajfEAl7K16LocWgw1WSivTFn95vgJoPWl3Ipx7VjG8qgQyrw4F6+ScwaugtMGr2Anc702rgWY
AyVnSyXFzWUyX274cEFeb9+4Urq7b6oC4ArEEhljeaBCstTKzb80ilhmMeohbnX2BxMw/BEQ2CF4
ZJCB5XjFpkVjGdONxa1Bf/L9kzUtvNJnjpggfGf6YEolBcp9x5zu+axt3dxaJVsZ06csEQWEs7Am
SyLwCdf77WeTl7/vkhYLVwVCPgwL4YZfOad6wfpQeiHAthHKSfbhJ4w97HkcMjr5Pj0NgBWVbXhT
f5Y4yMDWfj2UD4G3Qwl8DKtlbBfBhdc9kaB9Tyj0pRuskS8gm1iX5eCnTZBjJ6sZ68ZOSsCXfUJY
QTEMOGGkkHAXwB9zbiSBv9L+x29Mofbk2eWauhN6VgHZHpjgAI5+J//6s5+XJS78CL1Rjay/rb/H
Pw7zNFySl+jwF/3UhDB7Fhb/uclwjOuxgN9K1vDY7A/55K7jPWW98GUQh6ItBn2px9ieB2Kt/20O
P1G99QMQwf1AarC0chC3RnY+G/rDIIZKqmHRlJ8SyCHnY6grXbAI5APiCiTPbWvj0YGlf/xzwiUr
EfGxV+NicATiO+IR2YCiOQch9QUnnu7oQBLdgtMT0MhXIhwL9Kpto57lb6a76fAqv46okOrJBABU
jeaz2itqtD60KstAKuP7ZQjRkIvX433D54UfCT4NhrqFtMlau2fhMw3sk5mStN6TdTG5nmaRYGiE
9deJuZjx6yGM6ga9yAJmw43/ljnM1ESzN4H5kenD+2oj1mzho+IfzOLtI/zuzP5w/5VW+Kj8tBUO
nM89cho5ODD+VS7EdedubdJimTl6d5GzA4tYgWsrQNwHLQ61PMBCuPDEQ38Ll7ppBpp/olh90ouY
h0sUOfsD5wowuoj72m+hQVrz9PRGpFhDMWFXAvl7Z2WGzW6YqPkQ94uO6kRGyWJIPFmDppCZneIO
bE07kJ6MoHqof3ZnfSR5bzGvAiaiDXZN588O708q7ErBRc34Yvs7n4IDr8jS/OOW0wANhHNPLnp8
AIp1v9NI5g+SvdXxmizzBRrezFzinE1Oe0CQehbDDQ8qgOiNP//6SYEDMALYKC0J1M1qd/NgI2xy
hFIyh7QGTiY7bU8eqyX0q/yqKQu8zE4464RnIwDLcNp0CeLtNcZJ+7BYsYury31/iyBuzshlocrP
TMvfgWY3k6zoX6gaVUhkTKgMv9rEtDd9rJdHD2/EwnvPJRcfcFoY/ucQywBoRd2MV5r80AsxGApo
gd9rN61VaRRRi7bnCEXYmDomiV9lmRKFJCJ2MZLYusQcmVHEWmumLqCFo90uWRwQ2j63uxuMvwmY
6AVLmaIX5bFZUESpbe1t3jGYP7PoT3951noBMwuMmzhazL5O3rEBvw9wIDcusx5w7I76cJA+Bxg1
9OKAFT/4JRDJs10DbC8Uoc+myj4MIltnR6U9bvK5t8dG8jmV9WJoPUViw5z1sGuajikWLzKi/Ddo
XqMg1LmF8xy7wLdxHkG/8hD0mr2G0mJ+1En4Pol0Y2FzU1arhDMk7Df3Ldud0FX9mgJhPYy67ChT
uXcdoNbQwFkHpr3OhhyTUOXufUeWlebPdjsG/KRKkE6WIQMbbRJ72Rdt6MhOYzyptN+lfjRHLhrJ
rp5RkQG6Ba1EUPKgo9NDJsNJDmaeEFRA8y3Jt6IKlLHkjRdW6H7sAMkKfDoxQIJpmu77EC+whUWF
jIVj6adUBtww08Ktwgg6OZPo1Vjqw/dG6Li9R+Tj1cIul6A8HEmYCnYnYx1wUolISqNMxkOz7l8Y
vwVWv8ty7cNpVHvxPze2aoKeWsjpfzAqvACTsHzXhW0gUgiXDLBuAobTss4E7BsXm0tM9n4ku4q/
VYe6w/qFCOo3+4JtHhI9MrjQhZW5KLgEouT9f8gG74M85j+Q7zFNgRn4CFSUDznYocA9JavDAHxh
mbPaGVUw3y6mjUL6C7NgaxMnT6w8A5b8N5e/D7wQT8DM/7f3LwjHEank7Hq/e/pYK3R6N2tCB8zQ
eSToShVUuO9ag1pmQNz3wqwsBxs/oUpN93UQyFy0hLZfq6LtoxgFfZNm90feAngYb4PHqF1IybIL
fHUAi+ibo4Sz44e1S0O4VTnpnYj+ZN9TePahrAGvVEj4jXJ6c0OeUklMxQWwLMfFd0NDan1sOp6G
yz9C00vie+KX2A0yLNPbARRqV6tzRQAIK6vGDQOoE26ybFlYFn8xcHlDGd298ZGu2m8lpQB6fw78
YSvHo9+Jov0ahnlec0BfozfbsxaV6dUkqzSJjUaff9Luqn4o4wtvIkT5C1O0HL0HikmWMR+zt2JL
kpbpyp12GUavT1a6mQ2bLZV6XOUpUDOodKlJVwVFMWqEHbxdTKhssZXDL+SY5rybSzENPAk0ipq0
g1hBI5QoTU3Jo53hCnG6QKXlkAmW7NnZRnqTkmmuKTQWzLqMVisisf6hdbbQMEl4KlkQGcQ/CJjW
KJOcEKqz8mvk5+nu6zulOwoF6V6utEQVpxH4n5uWdhU0kLX7cZCdYyAgE293/3e+OwwuKiwV6J6q
wQ9fhCuWXKE8a2kneg/bWHBF0TwgQJC1Tbljz3l1Hl2QGW/B75f65s/v1dmCLE2zshDstRuJ0dEU
x+v7vNCNk5plnj4PCod70q4ndYCt37VVfDC6V/JgtkaRSbgaQKxHtR159ZCRvXl4rxq5C983qlyP
4zKHOWJCaBdlxI59mFoHXnjCpZUAGaZuPFdNBZE6ETnp+0obWEq3DW4AWtDwvhE4bdSWmdb6pegv
Jb6tazYTfUOYZIv0W9oS7s808CIxv1srCejsIqF1Vh3zCPyVwgeSYeePgozm0k0m6RVVjUsJcrU+
nnwh1WbuCx6zRzsdGaLOJnXqr2uJnX6ZyJJVFtI++TDlq52DIfTHe95KmzxBM16aMVnyQJx8KcJ5
a1sOYkyKKbF768XpZxYubOZOBekZwlmfE4lZQJBt1PQSULL0LlfOCZ5lvrWpVWl4cnA58yPUN5FC
idHB2fsIZDAKxSyzXqiUVDTH1z1f0NTPA1e4892SIZk+6WcsIJc7D0El8i0Urw09n26JEg1+2fkS
A97WK+IJzStOG0aHkY61AwPPz5FdWU3pyKLAHgWc02RsBKeAB2i1jsAa7SxZSd7h8QBhTbJNRaQx
ohJ6guSWPOQDH7z510urA++VfJEmPgZvTqaxGoQq4sj6+AYbaZR6YHKgtCEguIgimSoMe+8o8Nsn
pGbqbaNVm20aX44YmeyLbjSiAYeD6U99XZMKb6VSoqxyfoSgkK/fLDMI7+glOOqIW0R/pHKFPVj1
XDnmtlWiBk7ZTc1vPSL4jMddfvk+tHU3k/EYksEj12pqkH32gtGmprWrDPyEftWRjpaOip8eRN3o
RG+KiwAHfpRyzjiHE/LecsnF1JvMGP9VCP6vRjW4F7u/p+6FQ8Y2g+jFsjfcrdHj5D3SdEHk9+E8
KEWp/t6FEIPJ+1pX4R+alyZFIEohug0WfBtV9YmCFhsdvjilBP4Evf1B/FR4zft99VK+S0pbEqga
45kWryjlH3p+cHR/qAjRFy6NP3L4zrsI0QFh5fCjaYggntjJe71FnMuPSvfmMSTm23E+Xml1XYBN
of1RDGmQK9RzIjCAGxOkf7yjpLwaFu1K4Vao4Mdz6D32HbeQU5O4FrMi+N5kRkg+rzF81gGpgf93
pRLZT6HDvhP8MvyUB0FH9NcEQfsR5EnDnthAIhP23qSTzsELvuVnvsgLllK+AfzriS0Wm1rowJqU
Y9L5FFQBs6uxvLrowcud4subTo8HN3n19nj78HW0sKFNiZx6QEIguek/I+0oVHnPh0RWO3vqwBL6
CEW117aeIoykiZMSw6ex+Of8Hp4kgGjmGnImfMks04A5+Dom63Xhz2qLeuRPJ9s2LxZ41W1Vo/rF
QEDCm+t43o1YQfbDvuHNhFr+2a0L8p9UcIUjUV1+GQtTDjXmDHjVlqGxUfb6/Sqgatxur0Pfa9ee
DGX03BxcvAWsMFw84Nt2qfBP/ISSJrCaeOp7FA4+lb/SXZi5DdYYOezeRetcYmTa8GxCt1sZjMBw
vmfwn6DMMW/ujmVOhDJF5dTElWn75qTY/Vss0zsT/p0xdEB19Rqn1/UlseBwXQmzcVShNpo9GFI2
bUY0gUlL7kfdIosum0u7BftrzmquH3HSc99vUpKgIj0VovLL/kwA9xOioVrkU8cOWsF1/RUhA/Db
tJUAujaC1OhJEP2FMBwM/1UFF9jqPGpPWkyGbivBKpAR94wjvuhZZ1GIS6mRM0YA8BgzqfLN198h
UNMDIMOPlO5utQLi6/CbeC1yGSDKXBBDp5OAFkZ2d2jQaMjBMEadbnYjt3YPCmdeoVB1r1WZBHjQ
/qQEes+FnCi92VaI/C5KkHJ3cC1Ot23mZw3IBHbaci1o+Xnn7NXrElLQXs+SoiG1cPq/D7yQTyPU
Y9HsCiV7BX/UcRO2K2hizNECtmDWJNpTBZEm6SDjGszHbHYmXuTFf78xI4uETx9BDK4nauILhWHl
8QUEBiit4/qOnuioa9zFI7rFLcfmBztqXpG1BCBmK1MmVdj4UPlSjSzr/pyNMop0/i6jQv2HOH/w
y2cObu7gcafFjS7CeMQODv9bcVFpt9hMbfMiNowAFbAKnzSksYpbOU2o8w8/fprO3kxj43KgGv+f
Wa8gjirKrWEKZQFkfQSyRPRLcKVbHo0Ds59ibE6kbN0PLFVtHd6BV5DV3NGYfSeEiV8H9MI4nnya
X3gw0OMcLrqkpH/5sQ514t0+50rL/cjNb18CHDfiXwlyiaKvGM594yayZW4eFsxh2cZ4EXr4++Zn
kqFL3r/vk1qOysw296wqaf0QUVL5SGCX1Z7yso2RdiMrXKpDuuQDKEBjVRvUFwnsHmdN84tofARH
P2We+SY7vY/V2Eo6eDhWUSRViXSqCFg6ODPVHTLEB9lzBDDX6OFs1U+ic9Uab0YaGauU8QJd9M5Y
sWLF/LYNx5x8BL0X034UiqmlbLPVCm9NLb607sSZWHP3LzVNx8BuAHgobrA1uzwsblSecPs8ELJB
G19nkDYDFD1dV188uStRN4qNg0GZ2eC7IT87I6roB76MpOqitpfl7bnQyTYqUigY7mEnqVaQOyxn
wMAELTn9cRe/M70r7C8Uu+Cnhi3D9iFQoj4oIH83Aum1anwS/elQEs2iNf/USGtKDFAIP9vmA7E6
amUUvs9BPVBAjMA6Hg/R/xYNkOCQpm6miAiN3urJhCaWxDcZMzOp0k7VrsEAW88L7nFL0ks4D+IJ
v6Awv1pfGE1OqRSc2+mmj/yAmAgAs2VX3wEUdIpolkCyVG+J2bPQZsuWHf7CckyQtlu8xfML56+i
Y/T6ZgcyX/zZBxrpS93ZWy6VXKmq0rExdDGVYpsRWLOyeRSf+2OOu6EG/bWGVp36XYLv+Zo+ZaEW
GGFU4uiG4B4Olb19L0BnKedTT9n80kY5+DCgdoe18dkAYKe2Gmf1L6Mfh7TSgQfpRarLOZ1Nl5Pp
YB3UIr8fny4IIv1wyrQHyodCSo3wqs0EhF5MH3cqJp3ITHX7G/zpPYDznSEAqmyuyJYBt+QxrXRA
gQRVasyd9lJzRezmGYbzSMBpFbThuFCymSlq/hoWPKwDfZGyVLQQJFzDK6EAnSJ+J+qykyCZHD+0
9rA/pvbbILG2AQdrWuUoi55qAvtmgPS836W11+CK0j17xMfmCXD0vvV19/uCJRjgAG9nRbldOK+C
adhbiVaVYwytM5vXvBVjmb3gyFNonHXHDv+YiwMradvYBwUAp8AkeewLnIFdWpPUkjc0XM1CFzOj
AMKCXSz1H/xkNj2vN6P5mMd+cE9S21elZImBrXZ2eVzFikErzrum/P6ZuWE1kzlxm3x/2OGsV9AY
YySn25Gc82+/6vbbpxKkocpN7J9MZ6wMSrAFj2EYO5T2dRHZWGf24wtguHo3RXLCNh7RU8oAegNh
b5krinf74BRdhNk37j/zRPRs3VpomNGHrz7liii65NRL85gymzuRrV93+pauKX0gkgD+W1bJMQoc
S5jsnRgS30ppcSlpm2cyRh+taudsUsv6dmWhCMju4QoxDE0qunCgu1CpHW//yWA9g0CtJM1PJOJ9
2cfCq/yrBVO14h+CT/3IkqOn4vvSW0tp389TXX+zS9+PeLxZg2EiAC9bY0AiHStcx9WNq48Hz4qu
E4hVEi0SxojGe38mYsIohRDQXedQpjWRqanT1NcZXS8wIIDevXoPqqi1Yv8lR82WsieasZ187ySJ
tzHjiJsD2KeL6n7NChfB+om3/7QuyXpGQBG6LlbT2REvB+/NK73+XpC/9azpWxlng9AGqtiHRbnG
qKvT5axlSA7g5MyvImtP38Udv6Cx3+RTMO3BA+DSceGk93krkqsDhugYQ3GmfV1USqfGC98YCNZ7
KZEyEK8sUw54yULsemvcPOhqibkwtzfcZ4qEyZ2qNILXoBkIlNdyQPmXtzaYqIXex6bNkopKu9m3
lF88I2hJL8EtOTLER5Utn1D+J40zYWxzCC+RVV3QiK6dfamLNLNSVF6TffTz1l207hXi5UXpUIrn
KusoT+v+1+Gr37wkZxc4WrJ9q698BCRYGwrzrWs57LtWFjEfEXPvmd5dflLcbQXM4IxQh9tZ4juU
+Z2n+9CMOvRiSg2i3fHv1uoS//OIqPO5xElpQ9o3Pzm+1Zerj/maIx3k+F05/cLPEiG0VpHtd4fy
ZUObBYKrpsVXfp3+aUft1SnW8M/hBRNUVqBDpTKS2l7CKZFJd6h48eHEuPANte+J/HJp9N+rjc6w
yNlAr8H7pG40ZMFWAckB8Hef+eT4GcPY3Q7LH59J0NgN5JAA+HO9APg/WAOQ4H/pAsiUbrHApM0v
spuDmEOH59+jq17E6vySrfwdgEJ/dNAj817BztOSju/M0OFnOS/hxMKqkm6GJxodP4mqAxRSn9Ot
HC59KlZtvrnERe3Q11utdjIhlrP08mv+P3cmScJrfKcFIjuGuVsmErS4uqcNUXoZSJELGBdtDaoK
54WwT4AhWenFuRn3z+YUyhNpa30X+IPVQOtFmRUXrgHHlVt77o4tNmglrhipMyhlpUChCvw0grai
AX//90accPCPfvo4Nz31vNGELE2TOvH6x/er5kpnk8hl8wwDTBU6HfFoXtcevJJm1faFjwIpaQn1
D0OuTGOd97z0CmNv8S8AnZlk4BShHnnxZaGigP/y+q7v503U3OTubcQSLQxoVMBoq+qXDI8HLPJg
sk9oQMK3/muHhvzYlnpqXeKxjqj9f0RzpYdtMqHEeh/5XXKCJzeZE6zhX0scjOvDRBoHTuU+eBs7
EwmYrwLlwO08kquljbKjCJYfFRQUPhroLBL/i8CJa8JUIZtgTYIaZsegsJ3kieLK/pkA71inCSzE
LEND7TR8VXHLQq/bHGS5qsiyC0RjcdAOaTiGbluQhxW1dmQdn0SD+Y6vxMxTvwCUid5BlQF1hDv2
iORRcROMCDuAUE9GwTJE+G9k+fuFNjfHTFSt8C/EQ2WzGWWilWszcAym+7yGZQsyR4HnP9G4GEjK
7FfFRe7OiyTm17tjlubjqUOmvQ7zFEtgg3gLAnn4kYRjR9ix9O2kkDZLYsNq8in0ngGP4CcV8dsS
Lu84aio9Q0tiO5tnlOzfIQrkPYFCAkikHHlkuLT+fq0Sn0KTpBhi7Htg3i1IWe5RYHAQTj+6qoqx
j5o6DhTUuBrfcl4+tVbzpZ+nEH+tzTE1iIgLGNi8JshV+TZ2xWQ6DL4G8/GwDlIbtmmTX6oQPiEv
7Jfy5GsmN/CCD1IJDbRRhjP/SpgoIwW8HS6eb3T5UrxUF5fUyM8qvwx6wFB8zAtgKFaEQqRcGpdT
58yf99hVjkEJzppD7s+yGsMT6wgv00iLG0jkmNrGMd1k3PpfFYAVvHuPeKESPDRrNZf/oHhPpdKc
kBvloAIiy8J1fWYurB4D9e+NmDhRwFWuaJB91kdZuS1JvJFxWAcXYxTfGVgS4/DOPCo8ASEJlDwY
Ys/krmyW46VSNCe5sYKY48Uabn1Q+RW8B9jBq9eFtTQiBw0ZGI2NWph09P3H7msA2h5/AMS2WXq7
pPFtuDrIj0UrxusXxkWHeOstdtXGsMMvglA4XbPKaF5jjumko5K/GitFswgWU4vA5dunPnwlY3kD
cQBa64QX3EcP7Ucr9BJPhudAo5OhM4gkjAUSAz0E0YxivrfQZOdkaHAWn3JS3HsJwMRxGi6qpgbm
Rt7BpLLlLgycqCS5V+coPXTz6kc7CxQ5gwdNHjPRiA5LJIQFW1jeXtMnWEPKkOHpgy+Le6Th5brh
85sLrKSYQCrkTLab4ZHWtgblgzJ20qxEqVL85MGkaJt8oPyFq8Jb/UW+oxr2MyRLlo/+igZpGe/r
PWmPizZDqJ0g84ZB0vQcO0fyJPLb9Q/at8gPJeG14GLfQE7fMX5VsL+siV7TOYQzddDvGSa6x82M
4luuDnZTfMia4gzncJz1Kj2y+VmkpogkURgzXD0GAV7R/Svz0NkLYpkyXHWFONeIc5DyCOYrP9jT
qjtw91A5AOrizkdQ7N5ZaVPrsVUwTP8DTL8VtLtLAcMF0Uf/DGmTHwKdzuF9gxQa2jW1wmIfvXFq
JXZ2P8hCM27N0TqaKnpGar0PbLgAS3tuKRmMe1SlgY99u5VikXRx0RcrCw+dC27qaRlj1txSFUMk
60oIylrL6e2VAOOE+GIhjRjXiYbd/44YSU9qo7xo8EbGq437DTEEQSPoxLMCG+sjAXLhc9TnHtsr
tZPLYvUwY59Kz4iM8jb0Ejpgm5IoBIPVQrqLAn5ePcFYIcpsjYPke6zNmbqIm4gt8E7Iyy0y5sjM
4d3dRUIZu2/J4ANNuqiBCt4y5rNosbDvCASI5FGlE669xyK+euMEBAPICraSxw+JIRwvwan3qG87
ljmz++T9fRkYO6ewdzNEXzw4iCY0x9qvU7R1pncajXQhgdEl4mZQtU+yn1akfw5poii2kRBBCf8M
YplYda8iqkGc2A+V+NjHv4UyYCBn8YClmcWF0bmlklNzxZhnaKWDd/WfZVWRWGQnIC0X+tjj+o2/
Cul5Wqh/4i7MC/me/wL1QmcjLexdmjV4rSMgKNbazGT21Sybj6ry2FDSRcZvKtAZR5/CNeGshn4G
nDzNgUfC3oFrY6ns7rRrWJuAT9BGWdscsRxuGBGatvIDQbSUH/DC3FaXMvMd9FXRiAFLjlYKZres
w4iVvv5+D8RbBo5JxM3qZ/5wbDPuG92k66tWHxGozgPkrn+JirYBsiMCdm9VsDO3Lwc2Y74mXEzs
PN3uMsgsWWJRDqOJXsEDwwKo8IOKUb+RQA4Fft0xtdDgaWNBgVgSGxCN4L4ojTFxgS6NVCUqAqJ+
X0kkZqMReivqOk51558cvNsf3iyXDR3RtJeGoQ3bkdNinfKCrhNjvN8oBqrMlrkjlygww/uxa4SE
V47Zb4CrIiY3Pnf5D/9tL/wU9OKXerTzv5EHSfi9GdOV1n4DUD1PaiSFpBHDb1uhQvMXjAgeD9/9
+UDuKuF+ZoMrYxS9jqc3UMJXGZ4lW3s65PceCGapXj5dIABIu9UooIZUJmw+NnK7LvTYS6ORo2JA
HD0sGSxpPuRPMWXGi5ORbRPyyQPGAYAuNLA/LJIhzhHJTUOQ1orzPhnJdHy8I5F4DpB5UTbU6XcJ
GrcCr3F8Z47CYevBiqGQfMRI3lxOfxKaEKV4s6e/D4MiR8uSxN+7hgJUVvj3lsEvdbkiE349oaH4
8KAJDBqihH1RelM/39dM6CDhWFVzTjKuaU8jU+dDwFafNJxepZ9pzvkJtrJwb1qtSWBF4t//jjHi
lwIH+ICRz+hBVBVn18oJSKAluP1Gncqic1+b6H9mXqfcIQ7fKGAA2cb++2A8XUP4Az6hkFJr26m2
DNc6FhOpgn1cd9K3gY55KI7da2/10AKCww0zlV8aqhnc5ZyrJuWxQqf0XmwUjM+5sK8SvhCMx1HQ
BmVcgaAJvPZQb3h5Rjsveyt2jNAYCmDiMg2NkeY0xsUBhr4eUqrt3Pb4+91Csxy2qtC6faugR0LR
TkI2FdZxQOYXBvpmaAHc7XpaTjNDv0kK8DOnngLxyVgJUuMtShHMEFOqLhYxeSlPSjEAYEKNR+wu
ZA/aBVuYHwLZb2VtMnFocN5EEismQ+NRpmfdlhgb5b0myVXga56X2Y+SFxQ1n2guz9lwdJD744dQ
4JXDBiZUsqqG8u662GFMjP9DAtgi6l4AaqMnyM4rd8HUbccZO2DL47lOeipq07r1QMP0w9jItkUx
MjD+pqf+NKoFFKw7nLuSLtVZFcOzhZgVmEcwXJFeefcTHF29Ds7wTbiXlU2oISCV2k1gK9dczP7R
P98cnaFz7l0wvSkUT+MkeI6UZyCYcHlVPHU51K9wISUgnP4Z7a5Cw7rOyCiga8Sgfpq1dtidxLTu
aZfeMC8QAKoAaNSXt3pbVfWe6VgNqyfAarNspLfeGlLakz923gKroOE7bVk42X5gZWtYCZrIAXuI
tQftwjZjoqOEY8ykE2GzH1hRQ/R0nxnTgsgbjboZ34UPz5qOI2kPfjvzSMyG9C26fxI4+0Fcr7rI
+BaJK6riYenabG1/JnjyUTozTtzJM3Sk6MMkynC59jJKLRlD76zKzcfuhq/4AxRC5qjgVRNFjcKv
HHYWBm8RXEzsfgp4gOsANLr8e4SLIYGtLVV4ZmWnyU+qnQpKOrDoVOyPJAqwvtt4dRxfc2SmqAic
xvhy2UC+U3w3600/jAqGI2fBuO1SI3TJ5nreZOSqTffzVXonLk1s3RFRpMARo2Jcp0BdSQOyHoS8
tC0hmOO5wgv0kgt7kFEF0meNjqTstOYfVGE82/47P5Hlo7RFsSBYUP62yU3uRm5GnBSBhDt+Mpv5
G8zD1T0BXvFfvsTRCyvBONaqNwileJMq46dQET34NG/+DNEXTPQ0ADTttU6bUvTtLzBomBxTwUPg
C/uXVSHQ5b+Ij6M1mGGhOIWSrptElx/gTvDjThF8Q9VLrjMAgKeMuXVhtf+1YlyJKeOVqjiahMHF
fgWL3sILEgH8IUxcUme3ZXeonjR8c0MRlCe/jMnnMfPR8HN1iipnU1wWLm/HMghCisNO/SPKUpPj
u0BJUIL8RMxWV+yzG2RZ3UuXTlhVtYwbYKBP0/8UIfv6y5uGNqkQzROBPSTYavxFvefjPbTriZtk
wkNIS+mesU+sVlx3sK2h3dsWTkOxRXDauH083VMsq3WgzDjta2IV0TrgyuYI9sgJfczLVv2rbqbA
Ga9yMglzKqxyH/nMOwvYF1kVvvgXKrq7lPsky6AviD8ZLvxJACOosop30YptIezdKbLnK0hfkHjC
xqXp88mt6Hl3mAhVCcU/XKzxRzVknhyMoVPevw9V1Yaa1CR0qLevmh2LTZ9519ipZmp1Ve0UDyFz
I7u5zBSxmGK8/2G27aLnpUoSO2srX3w/g++qU1DbqVDib9vi0kii0+Mh17g+Bv7ac/hzdtR8gfPU
kyE/qfTVYhAOwSGmFuxmpoMxoaKYy/0Nlr+cfjQcYPF0dRd8ShUdZVInoFxg+LnrLU6k3MWVXaE6
FD/YGilgNF9N/P94PUMpeVkB02L+8jF6ONBVrIV1IrBy+HeOaQnljmgYBL2GsslRnRG/7vKFtTJ3
OehbiBJGjdlafdL/jfSAgN42QURax1Shh5D69s/RL/JYDqNSe4FNLNVbhjkoCmnS49qWVkCK/SQS
xee+ANOSnjvZGW3udVJTPaGeSkiFPzhx9Z+jArqgqjyHyCZ/MmQl82Eag2CyqbvWJiOWH9AG7u3j
0n/r5w3Iod0JOJbHuoK8CMLg3VJJsIqbgqRasYsg07CichcIIiHwTplP+PUFL2CccM6Yt0KR0SIh
QQz/tUNpE0nZ79N5ddLSfR7LIpbKXaT9Cd56E82fwaqy1qrb/QoF4xLxoISPtmqIBwozvXwN7Cro
Y+fUmEak4SeJiR3EzlJFcJP9839nId6LOwpBcmAOztWhUfXhBcUXtyU6v6lTpjbpuP1+xjRZ/h1v
y3S1vzZjInSlusWpEE6dw6oNe/Qt0kuPHWCjOev2AyNt/mMDKOExYHODemOuOEyaa1rayww1aoB8
Lw49dWoNcIAfXOCpDSqUCBl5jsVpjfqNvR0bUdnpZ8UkPSjNhJH5LzTvSQTXBF+KkIMGNz6VfdSZ
2KpOo49levA1BXqcVNVv0MGPPfgHv7qAxNwHKeRGtT9BvEqoaV/eoaHcKHERrAKjCg00HY9uD6V/
ZjTbfgPWaE7dB+7MPq9gbdt0QwSwB/qerVngxRUxbI46E7j5cEoLFc17hyfwaErwgQ3B1VGOQP6d
rNZIlpS+fPByIofIokUVD0GzKPk4aJTkj+97ABaVyMonFs4TMuWZ95sqm8+okX8Y5zcmXSa6u3zG
dwVmGHAE1aIFO7Bo+WHONKVKFSC6tzc6l9EMaJ8flEpZMehwtX/LuQ6WavfdqUanYrhJmWQbnd7P
iOXdQQtl0jTrX6Gz5mn9ONvebbzdivJH7oHLjleJCmGWr0Vaj9H8LDEoplBpgPrhSylSCHc9/1He
i5UAlBfWkI+6kyWePj2NIiqE+ovy5WhQiK/IhKgU4W5Std9hGTfGuTqwwwXlLs7pfnN7tdQn6a6v
ScSI8BnaJs9dyNYxotK3Ng37pS8qth+HGOWabfm38HmaCqc2tYXsIxkCzewlexFOa4mBY0OIUOYP
p7L2th4UuG+UqxKJt7zubmTJr+CzBD30gKoMrRW/9CIxhKrb0wnqnMdI6KYm8mPagKildzWcPFAd
WeDWGKl91BSNiMBGgw6CmpNTqsG+D5YPTWGTlgs/DLFUct44SneN93In6kyywJjpPC4lqZQn5H/3
69Z74tQFKcq4xgruyJvkf5OD+4Mlz7gXn0PWYU3wIJCca0psvjfWX5040u9a6ItySx3BgSwuXRxP
R5HmgQSS9xE/BD11noN5Kst/My8jpn77lFl8vAPK2qXsl5Yba8xilUDsQqTUdEzGzmGTQ/6B0qvF
dPFYhItFo+wTtusLaQ4TkgIZ2wubZnkqDLZvGSfAyNGO+QaX8P5meRZ19X+AyDdmoj+airBIoK1I
EP8h/lgDto8slzRW7tkPR6MoFNW8ZETbZKat72W99KpzayMt6/yH5KzI397tPhrQAnwaZbyVoIgw
hlve1184f12MTsnuubklWRsBfS+2PKsRDEnepYpe16AsFzzdLRnR/ED5jpCQpQe7zmyrUTMyeI9s
GbfhNTBasns4Huxqd33Fas2y4oOxdDGnNzMli+OOaLI6dC8LtxnmBFhPddy7iTuQeVDwKpz4lr0x
pS9Smkb+pelbLIsC4XtlvZMJhmmIvc9DldwsKqiH1ozvff/8XGIglThRPm0uYmKlAqdklMZxFiDI
voW2F2jDcqj5GF5jNzzz+jzyLO3DnisT5BnY0cpDsAUgwLxyo7Qun4sk7gEHJUY32IZNaRrvZIwC
8Iqe1Fr/uBApfPLuF/3WZ94hLtGYdA/RcugGgYHC+JUGIded/3ii81nELPOXqmP6uuOMnr/CEtaH
2/qsI+McKKBZgfq8eJsoKjHhVIM6U/SeId0Tod2ri5x98yuck3+SHmE/h+6rjiPXXsbr56zBv4fu
LSSMa2/FxPTU0hSmfXy+efI0Q8duE+ZtrPRnEC2iA+0uB0dnhseD0yWOmMpzJTjou6xqbEd5mmTB
EloLQY765PT/o7QU0PYNwNaEEwbAeflrFVv0grXgPnDy5aX+uHpV3CISUENPzKvMPoiYqZXQnCk8
wv4OLjhZPFRQbNpejIsnjibS1PesveHnCL6T2Vh9SR9bBm99SBY8M5fxLkLy8wyCkMa1dMPBQKTq
RodCv8Uuq17wgwPmqPSQkC/Qxq5up8zqrZMsOU4qk1F4xZL4jQ0xOVaWhbI51fFUqCGlE7XeVPbH
PAwLpuKBjy0+0tsfMgCn2WYkS1R1Wu/qkm7B8YIR/osGH1V+XPJ3DmEaE/J/D2s+j7e+Hx/SiW2Z
3kDCqxWRDf67G+QUo/GBFC4PQzOWksMvLgwgx4l6XoqS/O4qWIILofX7AsDdjivLrAACnbJq+BLi
vD5zQoSyKo/zksBCTHSAAbMtTMT8rTZJMzldhKezyfwC8CeoSWgRNmyKwg132EWM3XA90TxSqAEX
F0MLrCo+hTo4LcmOMZzA+kAlcC0NqhaaNakVpNopR6fXjGc1XfVIyi72uzeJpLPcK851ZPyzIhd4
zVA8n53owFDpZAQiAlwR3agSNW6GRYumWhrXLq/dedkDawfSGWI+GUEk7YUowq1NHHAgojpFVt4n
xHDdz3e/JV4xI+6Y0vQ4JdN9ajTL96mglNMQZ4v8SKzgH6hGILlCHFO+toyLF7Zx9fM6UqAgoomT
PWDyXbIaYXcJpHS1b7J+gfnC/4g+6f6NRrlMtVkk0brUZhAicRNM2IEShFrLoAi6Ik4QQfcKLZ8P
nr/y4CpNJjwLvA40pSXrrkGPBKL4J1JHbeFuZ/Ra43aU3aGA1UPa5OgcZ68LtIocP9rIQMop0e0i
gdWvx7Kc88vdEWnatqcQo31ZYe1XLUyLIddmB0bRjg02G6UOhPmtcyPFvIxmRf46UUDKkAglFFpc
38xYzV5Sux5nfWoL1FLvecHFCIkmgLwsjPw3jKDsmqCSdKZc4b+2vLvSpi4XBkuj7nuUgaYG0zV5
nZjXw84sh1RkBZ8+6KNkfYl2gIX8DFfy8Jt1L94IKZcNLemAC81xobr3eSvHYpWwler40SNh347u
ZWnZ4Bee9Auvykq1k+fohwaI//Hydyywo3xYnF0jc3zLpw7QexUGSNe1uoyl55+VJbvtNEE51KaE
jxsDA2b4OoZkHtQdCjm9pagw/P1aBfAiqrm9+reaATatuE2PKn565+HD8P5jif5LKnU3KiKP4SzV
iQluIzoLJQFIVA2fPzma6RW24k+WGzJuOZowwdwFWjLRdDVXcjhNrW3HK7+Uo5EkBkd+we0o7vB2
RquCNSTIA2jXaiaYCwEbR3IyHATiNDn9ZHrnzI5FB00UDhvwSqnRZMVbzJHLrZ3TJdsgcfMhx8+v
NwkhzJTm4WLNj4NKKMc5ieMghRBe9OnYOvbKo4cnJSGOBOGzZrB8aG5RmTStbqqBwkGkZU2cA0zh
8HQW7DEvRFHpgfNPwouL6SD0Jn+MQ46PQbki59YCm8DGAcHTpy2nIXJYSswhHvk5vnE3dQXQRo8X
xBOUBO0JqL9paYzRnHf8qsnkaOOm10u3o7xTL0lYIORGzvCNBWBxBRGA/1mD2rqTnboMENjkE+C3
EO9lWxjEEmuxkg1RoLhn6NQS7D7A1UVSDMmDaQtWE339dN1UM/pAUjcszUiCDnD7URlqlp8vLOwz
rlUHkQ2wQObbch0fyfGCxnGRsp2LFMtEAA1GuiXXiTsLUieBE+Hswml6BFC3NaXveEoQzb7UB+4j
3NtTyH76vZdm/zEhET8AJQ+YFKOaaTV+Vi3fvyvawpN/Tl9weGU1nmfsC5ro+wDUV832cYBzuzZu
iTU7ion+2zA5BkZg0Eqoj1PN9vl1k5yHOph9JbsWLt1lttNQt6Lz/A57gnZ3g2Lty283d4oPKJRU
cB9a7LX5w4BYEP/trgLGcrW2OMj/+PUf8JFEhpTWmSAD8nO3rYK2LAXyubKCNUtVgjBrGjgpPSXg
SDeaVURIlFjH/np3ZQMdasQAUiYvQbyNay6SGQu01A/zzZU0dyW/ABSKRnsWHH5PFfgS9+ls3UC+
Xa6F7G4YP/3dnf8wJnD9wD8YFmIwk9T41hCtu4mZy+OIUYlRlIlrlq3+2/LzDxGMN8RyeWgm3pPX
74sM3Zcx4dhwbDV2BusRx9zIz7wPK/UZHejCnrp8uEL+25/DL5augg+DCSLbAjy26oF/d/kylusU
GD6mC3aivkaS3BqylNJl8JSfsvNhCaz5yyK840hVOjXOp9P4OaEJVBxPWPz96Sv71vNw4oP111f9
2QrVHs9Ra0ctnYS9P7KLW2A7iFfn02cUIUACHCTPhYVvLr/AC7AnnB7LYNF6rLcr3Bru1X3GBPGb
rr0PTerjoYQrNEj8rJGk/4c5neBfDDkOm7lwSBu9wn8oxFStxnZI6/yD2xZpoGKdAr+H5VJOP5My
H4dXQhVHkipHXfQe9uI1IHLgPHYrP7LGg7BV1jNDAkZp40tjn+k2rzYuVbXqy1xu2EivHlBusePn
d07ijkkzYfbqttqU2DvN99C7iTN4ocarlGYR6tfIfAyq4aOIwH5feOu3d6qxG97f0kSPzUNeC2fi
mZMwYAaEph9ngJAF3t+ciRgjD2Bwh0oSx2rwG1EdcJmlRJh6LdO87sDAc4fj2zwH0fCyvQ9H2stb
K3V8KG6BqtwxXNWl9U+d7NptvjPtrTpOvLfa/fZrlnhKOuYUuXt8qoXOcNfm8oClv3wnp0wG142g
FbBi2lkgFFoXbXShuiqbK3S2frPQWyAFvxbZMpdCg9OV/f8Qpof86SWhlDoDBpD392zXvCBPUp71
RkIljupjL3hEFbernA0CXHy8/AlWGpNurEk8Yz+3lyu1aUu3pzDeUBZENc9UEq55duXeX7dfLyst
RiNJKnd1xFhIoBmefhq2rING7HbUyn0FrWVivPOKdUG8nWDuGX/8uKr9T/gDDiWj/EBjZ81KYo+j
mn4nUOf6buAU/hxteHvdoAMIGx6235uOmeW8dIFKUbSP9cbuIOei1SPF5KfKXM8e7WeSLXSJtOlq
m8ez0FI2NhWWePGv5JNvbY3XX/db3fyDBJmNtT6k/kF1/7C/1L/4Z7FrTQP5Ojk9iGeYO0VmHYu5
ozF8mmfIOP7C1CZHgQyU820gstPOE6drvSOw5zS76UK0VNtZetK4rn/VB390sgUX4SFY583NpzQw
42tmDNX/lfg456TYDKtzLu3Rgaxu9N4d//ZI7LjonDbfjV3cPWNL9B8UVhcnSQqGS/tny0wmpe8x
SkYv2RAa+ZN81NWrFSRfThNjzaiX+QiCHAJzE/uBiMgqbBDoRPpO7/8P4Qx1LxUvAA7IKrIxJUJ0
RbZT167biB1Mdx2xpNKLykV3CUBizj6wvd/qX/TuzW43lHQ/uVmKXasD17gsQOiDTJ5j4VNGeIxB
R4MXmPAA2WBL2l3+E4jzlwS7bgeCBQoCLrBXQYBesdy+42N2f66TNPV+qBls1maoz6E05d/Q1ng9
0dKzDhHlpkJP0eUYxJmVb9ZPP6Ur1AySNawAjHYhhrD+LNXVAoBitGUg5Z66TKI+O6wA0zITippg
rnrBYRxS8Fp1pravxkzStNRk9pNdb97PIFeQB3K0bIuGN4dzcQPt0nzhEj4x+qYdRliH0szxxGgt
RArUJGHyeLEwEGz3v/xwBj7Ql2MdlJYPdn27aB9fZTMHcs2Fm274fOCiU7UFam7gzUPFDPLp5nLC
QUQSxoR5ng+3zGQJst6MF2SaCzEpvdU0ShYbWvA7X76vvCYpUTcEA3NZHYq7NDhaedy86W2ezwIc
UMjKDFnc64x4hlhNbH7ylOsLUsRtDbUJ8xV9hOjheZYfluwgE5NlXDpuFU38tOTg4ubT/ax9hPgS
/yg5N3PYgcqE13AhA8iDmL27gt0GPOudXtMsdtMbnvW0PXzNMRoY2m7/FkuRGJFU30rkbgNDnzUO
+isuGUxI10SJbn9TNZ8k90Y8N1SFO/t/BKBu7zpPuY/r5Ph/q9NtuNybJ1udmyqG07QFS0qtdSzR
Mi1a4xOldoYYrDrbhQ5jetMxDPI9lXcyciCv4PCUW6vRaRNKkJRdTHBU3+uTWPsCCYvFWv59dtcp
+kF2wmcMctwB/l92Ra3YzTcDZYF/dBk0Zmhl0hT+Wn4jzJlYNTz7XtyPhjbXdW5QQAthgzyxJ+l1
rhzHxisJ4Pu4JtmtARWYy8dTWw+VKYEc0knjNsLIJ4IIDHvpI/jEUogT5IMJCrC6dlcclLuLM6Ne
Lbkw3QdEtGT4I5FUpfgoiYzZ55jdEcUvUazMAWnjwMzSxNe4GLj1AxGV7XiRVct+UNZWDNMwQeYx
5hG+DGrEO/cwunk1YXMIodCXTXCI9J2LzHFpu6BTq2WQCN15i/bfHr4cRfZmdZgDfDeBYm0riFL3
1IHkmcFAGzV7IaNkObW0Wq4CaoKDBkKY/VEMtdbnYSkKnjm++joVOE3yJ1f7E+CodWBzMU2Yvcnf
hLC0/p5dv1JOnb3wfk2pS1ZsJgM1ecxI0AG1XcWmOEBSHjOTRmUIOTJ94J05sGdE+WvBvOC7cqUG
Tx/72/RuwTBGR7WDRldoOr0SOGXq63itsQGD7qunrOamuBU4uLD7izqY8/8dw5OKrtNORZtCQxoF
j9AiPPPzutUsQgHj4wumG5xZrkbYaQYMyFDttkisq/kuBi8lL505bPNLPxD6zGyCLCYKr4x8+Whp
DYaCft21vVSieRbZ8CVcrV46xNmzF8KeIJfY4ITFLgMuZc6Sr//SXrRHZa9RpXSomTosZMRuV3Of
Na0ixbxp6dwpKsA8rwlyynaqWYJsI2aDco8PefxWiFuJm13EN1V97WNGiIe8klLJ5FPPwThouS7M
KxO8lJhL0eS5rhJEfK0tHCI5CjmlRjRATME1DS6/NbKDTAd43DvUjhtFho82m2HwE0Na8mGgwF7z
QwWIp55ms9J7nTbuSu2chSdDSEWW1KNj4ivpPI4qLO9mXdqrPFHtdR2GLOluxWqa/vz6hHmf8yhY
FwGvBuuKdmFvgvILdvmw9F+ub6YOXE2vOVMFnf4HciVHwt1PhE5gwzvwdC/dpDJzIiOmug29PitL
eSYmb9XPLcZU8HcXwqtEidEGt6yG1vGAv7AvTDvtpkoNiT0LJGptE383daaKAnWlJPMqQ7OXYE62
VTMFn1CujtWjISbOCQaX9t4ZiE7KrsuMAiCqYf28iWMzgXG6aOydYzmkTACVzsPDLibcnekXyW3Y
8q59OW7rMpqwVhuQ6yRYaJuAJkFKiSSpa4rxD3GI2tlTFT7eb14NWWgbTSWd2Jcc6zQC3phMcLCn
egpyMV6hCrqkDL6/JfJaV/qvOfOP8UHwGVdjgk7uQ4TOK7nh/Iit/yyJGilwzK5aB1qphDlsqfFK
Z3r2M3AoWwHf5FuAHHApq+aO6zcsYZLyckkBTol1G9FZPP1pqYrOwSz3n93fPrVa6XhdVcaJHzgB
5XZyhlEsNP3EwMyzfzBzMWKEiHZoe9YHUBGxV2jAgX89osXpbMcFB+90e7ViBOfwWe1hbHXeWAIF
6AhEXOGvmzppYr9d1jn0mN8RZBNe3jIt2CqObOYKh6y67SVgeapdiqiwLqViRe4yOg/X/HbUHUR1
8BmeG6jwSxFbzFT27TSjROGMk2K6NLCe66nZsh0OjR7yD/bEh1SelEk3aEMkihDSHm8PPMeeeDrb
OR93a/H7zD4MAjYfN8veZlCMdV7u2z1lgC9U35fH4SCaZtdgYwTds184od7dcW9a7F9RiCpi+llC
C+IfCegx7b3zoR3vlfjk5N/SvR0rVIzbfXkLv+hUhYkW0vvWY1BKE+W3WjZJ2fFqlhuPAP4fBUtM
zkJNC3Ko2x7dXFA9KV7oSYqd78A9zHAEkcd/3AYN1mqbmD8LcdLcLL5EE/BuPMbbKiGKhGaJPxW3
ZQfKJdVj5tD436Kxcy1dCRMY37zJiIWW/IXAIv6IS0z+ioXXibN1E9I2jdMz6BtUawuWA3U5nAAV
pG9YD4M19xpsyrEnS6b7bp8FWg+1cU3+Vyh70bgNuUTJcE7nQiXuK7oL5xL+BCHfrL6ZGu6g8DWz
UtEUcd1mzUomK+jbt0BY4avHoc6RJIrJybWZeDP22j9n0ZBUhaa785up8rzd1F6JqPG+gdD8g5wU
DMRbbwS8fkR4GqOoagJZQQIzKEEpslmEcDpKVhLpA2NxV/hckmXQT5EVTqfLHuZX1SXcdP++YlBl
39+xFZxD4n9e8tIj/PiIarmOULlHn4GT5KQfdqOzjravbUWmGNIL+8oT+rxcfYgXDpQcZYLG4g/Y
A2exiLwYDElozZqMAqW/Jc+heVaUhTZHOKoTeqDnHpH807F8vmHWkHbKVmgv457oj81sRKRsgAi2
MVGwvmyp0gwFJIgsK6jV2g0BbYxn19PCnyMyh9Rk0iEZKuChnLzlpb2ha1ShzRLFovq6hBNMl96L
FibqtOvl2pg2G/fX7Xm4KhVK8Jbqo3agpHFEsOKhtwLLSEuGplEbswzsANCwCU1RfZnZOuD1OE6I
MmH9yQ7MozgciidNgdB+XPE5amI+azc3ezLDUJLNiocIcZZNCAVsdsffuh5P1Ue+Dv2nBGzHsG8f
r3LemXMt3+ogCqEz9FyJOUynieLVavABi+qi7SnHWtMJSfTsIyG8ZU47JlFssgaaKLf0uFrBJKPT
XMr1aee3RSNoOSZcem+9Us+2Fuu/2PZybbIg+GSi+l73OyKYmBl+X6XehDM0kgNki/TtsmRELoZM
LX5UmYTjbujceDSL1BsQ5nvMpjnhlHduFrx4i7cx8D5q6f/lnPY2ruU1h3K+h4rh/9oP3xZx35Yf
L3zXHQKuUWX0vEK4HbXIUJ5izz2wg83w6mJ7926gRikspvhcN1z4PLNtcPc5LD42ROHm979PSnUn
60uYFlDNPs3LNTnRY94XIU+CkQQQswQ7Z+gwo3uGCs+0YarALMyYO49J1I0cd8/f6vJcRwfuvTRL
1Go4Aengo3HfAnQWBatPvZ3oy2ndLAbd/cnfygxSuFbZNNLJoFmMA8UNqcEZQKe6GwQ1/XZ91N/P
5XMfYbyKkaVJa6jmwsVKi+6pQr6tDDFcdd9Wum1IHWKKQTbnryqoj8A6alw8tH/s4g+Td6J6g6Jq
hFmUJRSyZJlkon9dnwqNtGBuloYHvS7dzjHwPWRF4oVpLtAMTndc44C4kE9xQS5zmOUsPMt1xM2k
AiiQObGBOGlHVESG8ArsJcto9VG1YcQsx4wl7lA3EsWESlIMWkiB+o6D/9APL6NnC99uPN7Ad2FH
20SAhbcWEvVJknEn7j8sl6ZtPBvpHsldzw8296lU5cGMrZhQ8SR6Fwo+MtDroJ0aqm5+v1wBKhIA
iohwjR6joxNIHforMc7osab2Da6EvNk4IrTHkZOTTf4bzCXCh1geHVFyOoTzn31Wyxyhf+9Ch956
pYTEEFghzykq27k2+fl0xfKCJDuejs1H/alhGeaH2JOfr24njCMuVGu1E7tlKaEleP+g5cmHO4pX
DNDOrjZqgbClWxTbpX0UCSYyBoYkwvE/DjTtSYU8YUnp7mrLFTJ4RTx8e9lj9SnqnZY8Kft52XG8
HT97H7/PCxYV2OEwfXDBTqQoxrTy6OMakj+L1y3F5GW6VKHfiaqKtZ4DqBLyxGwmi6SJi70PCYLu
wTI0tp0tRN+AWR49hZEsy1SgVVRYaNHUHPLs1nkb+klIxbOeV0noL3ku5ndfQ+t+Hr8lT6KS+7Ot
mF6lZWo0IOkaPRWpwkyftbdEgnxid27gEer+CqLda76Ds2Wv62fl5Fk9CiYmcCTUnSBydFDn//t7
8EOUk0fVTILK3oGu80jqrILZDVeppSLD8e9vc86M/ModALWQ9yGd5U2Yu/llk3go3u/fjmXOIlWX
x83tuzJcZMdGZtlKjYCjI/4/wC1SVoYxUtHRMLTbHpmLjxmOg/30bMZLtIPhl9CxXAgB5M8AkrMk
yqDaqdavzpcdQ0ZSdAw9m4ZXKJXnCa+RDaLLnSF98HI46S7vGGHBjrPaqPkiC0rSyfgyH2VcsAw7
jvsgAC7HB5j8XcUlwdrLQFKMl3a4W7aNNjZ8joh15hJUgKvtE0jGC6+jrwWs4PRnVs78pN9a06Zn
qYNiNDH5ZiVMOmOnIKFTtNO0l1f1oARVpQ2D9G/nfVZ1WKQA4VKsEa9SsC+ZEz9Zgedt4Spvm8wI
Mxn85vRmTX8CR4xRkrRyRKAVLVYv5eJwRsrtmoGefpchtNX+qDxn0UYI47Gbn/bGH0vjulXBtMFO
Fo9TMrLZ1yZpQXyRrF7kOZLAGPINSyjYcVDByX8fh8DjRb1xajUKntQJwJ+EMncU0douOcmZZPLf
PdbGZDg7adARQXhXeanJWvl5I7ytG6lfs6gg+9nHKllXZhumHYwxWrloS+n6hZoM3ZPHVxZzJTRO
C7PYOha+tnbdWyg+UyOknXHoelt+QxSwvfxAA7mdQbXuegawEOM6TDvQR8+mlyGfK14L6KDvf6bB
kFvYGRfNPeNHufbDaLukJeXt6lCTbz3GpIINZttQWkaPmhiDL1iCIPT7DVW8OS7e7bishGLHyc8Z
N5XtaNPwm+Ys3hvzY4ccutiecdW3u3bL4Kl5xqLmxHlcUvPPCCROFAqkunGoK+rtyOGF3eZEGgqP
A/bk3YJxRyUq2VaOMhjp3YYOeqwYyfFICOTXJbGRoRFEG8W+YI+2iVaVDgAWSzs4FVmS25UN+Kxb
dw6jp5zeGYLQgaeRWlVmCfYo4+REyHr1GCh5aDuN7OTGqZb3s3YAdP7PsxgOcx4mKPmwI+cT9vcE
xczrTvztiiSVubSSDb91tSU+6E4ldUmOagG2evica/1Nzc4BHoXXLJDxXlKh4mJBH1fSjUHZqA6Q
SRSFNBp6t6DTqbkGRdw0Qz5nAAb6NMcJZCz655DmYzvi5aaeV0k6xr/krje5phx5qi/cdCqn31bm
tTw5AYYOXe+wu/C4fWUTfGziY4cw5b9CVFSD83yIO1MaO3NRSquY4P6vrvUaAOQVHOUEKe40UlRF
JvyxCNjlXc1f2aEdhgRLL8EuS7SEu9HLByG7i8wT7N7o/O9eU8zxglN5pBoKOcPtsbe+qxvFJ48K
veMFBhdaPAJ1aOnEOhJyEkHIegWoClKv/qACoyIUoaA2CsUJSDbS52tqeYl9UUDmhNz4/cEKsskd
uRcs9Dk65vWT+Cg49DE9XjvLuw8Ow1ADdH0+ZvDaxx2k6gxIPZCWRdqJ3t+szvLdjn1bM1cjXWol
ybg6BhE8bsntPPuq50odO8uZjaVUF+c73RAX4trdt/pttsOujIS6LF0Vaey4SS07n+kodM8+yMC+
7wLlYJmKk9SzAbXRa0mlmVhz8KJk1k7ab534EA+fkjjZKqF3Dh3+2cXhzARbD2qVmL3izOKZc+1J
e6ZWPh3218HJyqGTLXY2+owVK6a3+KILLeBz/hI+Texfzf2PrxBM7qtRMqCYFNIJomPKS7QS2YsQ
DlBHmxkMzJfIhbiXbVBGekpJCe+xyqh2LMhgnCVH+tLoOCkujnzVc2SO3K8vzTghrMRwcHCl+nrT
2rQRmsuMy/q9kFonE3FoacFeGsDxMNcZ2ZlOAS6TU0GhX7eSU00HCbOQJzDSUiT2qmwc9bpXhMx9
CX/AS2KrzfooVpKtEQh2z73WboWgiFxPf1GoPd0UtuDjwb2Z6qEJmCp364A5cwloXhomAzt/68Lz
VdXd95rc3a86bG279pKY+Mexa0kKrlBbG5Drdx1vVP/eQacVtjuFukDyEUUXjnwPYEsoqv9UH1/d
6G7GVxkW7yFUF33Z/BiXlNSODTMjZzTQ2ABUmiVljPWX202M/FQY4XeDTaUPpb2m0MRP8Y5S1nFL
ISl24tNyXY09wafTGhrpyYWaSQfu/Cpgl34sjmUsMKXi35P6LCPw3L0yyWCjfnJOZHpT+721N1y0
VxXybkW2fqX6MMrBWDbIcPvIQ7tENSrCP/lbkmM46pQr2yk3XN3aD5kOXhXl9HArKriDoGCu6yoz
NLx6vyDirKq0aIilNwn97ci+c2019MZqIVN7QoFS5dDZ84KfLFHGm6QlLPa2XugW8S2SQenar4i6
OZWR5FA0CREEHute7uctHXYP1oDlh/Of2qGTIaNDPKlA3l4Vuude0V8gY5BxQ4bw6tkAYy0JRERk
ROB3vFJ/G8plLCo9TeQKuJuKpzficW/Y0C0FrH37GAfq+y9PhkICQWQPyg4DdJm3Jx0HjHoe8O3g
loTUnRZbdCPB4j8U4VWcrMJwqBIY3N8cOScpq5W2KdmWpj/33zc9DqyjVt8dNAPDSbt5o9RXDg1v
8IPsiBZS6E5zm9Wl9f5iBexkTEzEwn3eYrEJ++lqK9pIDgWvTiBNRdmT2S1Q+QwoJe0bd43y3oID
sILvtqZs5IJhaoCReg6EQSgPDgpBpm3s/ccfVKGkltIqrksC0X0WmPYmXXpHlZsUcluNuONNzJnH
0rUA5fe5oKdrRPIcV8k34QtI7QIbgYr5b+q74bDEaW4YUH4hPgBnCns7mLsm6C5V9V03AriR1v1H
z8z45JsqX0WoJAsMLZQtvxFClc0QlOtHj39FQxy9FIaAdsLiC5NH0x75HBEN2dhJEMMcCxeQf/QV
Urnve0kMMENcg20RKxmTz4ZmNadVmtP/XNM2kuUW0LE5yPsjLmZrMxQi3xozIX4tqQBoGKhGL88P
Zk89cUeHgXfY4c4uiNeB/oWW5lJYct/Qan18QSmsAtOhMqjPN7vsd2sAXSnY0Fh0Xwb9mJWqqxHl
evi0v1z31m1qkhAnxXbgivBUiT8NTOsgBGcSfScneoKma7VFN2ygY2lu8R1mwvLob/R7TaIbmE2e
AvltW6uTEcXWe+4xQm8rxTJBrXV7SJJjSZKDLFRLB3IGE1B7j7LgRLp1gDRSytvZXWAd0t5IdcVS
pu00P4drS6qmgw0ohJKImDjSq5xeUWmxphXTbh/6NEpDMIM/6ut3eE+nbuCyNh23BgsxLXXxUVJI
oJWiPsBi4Vi04s+E6Gn3GStMhqq0lY6PNRBbbVWZt1JN4Axw4KQr+VqTiTp4XvwMoTSC88qJsIA/
vfRVfgiEKfF6S9xU9iwfwoOtA6Lnsam1Mf0PC3Daak6WFGwER3vfzGh0Ln5JQv9z7oepBU+JJDS3
q0klK/wWJ4HGCOfn9fR1my8HiIADTypsx3x8TjMCqkRlfFQBsEWDTrH1syU1AhoixgKjsEM2FbSA
lsEIhTWl2p+b7TIeEKKybjl0b2DuRgSb1QG/5KxK5yROLCuwYRgPnzTlEA7tORsQK9rGQaDLpUJc
beaWm+l4RKDDH4o3/tU97ypdi+wrNXxcA5YirRcRUAe+Gr4NeQJAdzC8fXGfCi02qjyJmxUbgPBe
q9M/kxv9yG7LwQc5y5qGoOJLQu8XlCcWPsPC0pB0OWuabreCgrTFqu1cXQfEhrzMwOVvkgx2xCh1
MWfFtfrZXNCVOHCnfWBIkAxsCpzVxGql0UJqfBpjT7OXc8a9y2AXnNhHBXc+o23tKkD89kp/jj/C
yHhbuULh8t4kjdgdQ0WvwzM5UzJLq7AJfYYL4u0J3F0+6hwLda0C9Xp44/k3LFUAMwzPGbQ28gNL
+P5YbFGHBOkfkaU4WLGxk8IMVwIkBOg+yOy/E1o5ZjHjWAQ5w6X5pYr7/O9lTexpcy7Rgc121M9C
cVBPoXV6u/dEEaZ7Bmsbjnx3psIzdqLHWupos50ZNd18IYc9wl5ibl4BvPjwRXMqf46qnSJyNpH7
+lIY39E9uxe9myxYoAM2/lzPdAux+fH9L4CyHIBPV+njtmhOeY7OdVFn6DYPN0IQfVIHOgLRitkB
MFH33mW7KNlca3Dksf4H1S35s2xBqTnMKMoksBFjEr2Js+3MUWLWQMLO57j9SRW2q/XY+fsD+hvD
THZKKpEs9as9rxuVxmgcE4DMvhQdaeVc5w0iglt7tS/MBakmN5ICvnmgbhEDn39efwvQon+wuKon
MjwjbHvW9uhXL/9hbRVztGDSEFhIJs2t60QtJLx3/W7b/JohJBkD2Qrbsw3t6POpkd8EfJgC73Dg
0anWf/jDNnstASdGg09H1FJzeL9tPM8UQqOz80ykbJg4q8OHDvYJP3FKLt/+SGZ7UWv7/oIHanag
P18jukbelsP/BPF4Ss5xPAwFZC64f1x/NAXAKqr32Jr/UHvlEZgnqTEFGPKIXMneQIWtABuE5Vh1
iihESJYEy+OwvcWe84HOWuMmnPu82iN/e4Vm+S5zXaxva7LLdb3fA078JYj8GxSUvHADCst0U4Fk
EpRLOuYZzo2hq2AuJ987X8QwEfmdfvL9tz+1uSV/2+Wxa9KxmaRA6k69NVOSzZx9j/pO1YU6+n1K
31Wr9RgmbcSpFD5qwspmsq3ejc1UlmfuHEv7FlnJH8o+6xVME7rWHCvs4GaAjqxKPaZnviOOW6U9
xIWcjRg20wfYK++j3BXoehUQnmTsaG/0SFblaAMcogj2ObvcqF9rH8kgqLWMQxiHmlnzFB1aQABL
F55Tmprv2WJvDfyHUrtoDQntfZZUXF6q/7ieGnLB82+EIWQfxJE1VfLFZ+EJN77xjMhYd6mNYo2z
xcJpuqsMPoa1c+mnjH20lwVoYoGq+DWrs6IrF45QIBXRilbz/5tb44x4/ylu3NX4axuVtl+C579R
z+PTzn4TpQJ6eiFnk1e/9x5bdPnfTa2hs+71TSe8ipcpDKGu0Z7byPYqLzBisJ6ASncph/73U0T9
hf14bl0ZqwDzMpBZOPTEWOzW+6yTjnpDmKNQdf1toh0N44NLdEbe9lrvxoZVB9ctwY0EfzNaKsCu
XxCbh+622yNT7pGqNI9MCzwuJOw2Ppl2OBAPw0yZXzpaYEZ7/ts6/Y+AcsgYo5tbN1XO6vRbIWYN
om3WXlw2fEOHBCOW1MDKOY4AlYERgzv893HHypejraKTcshE+z6q3nwOPkSoif5GgTcycHBjx4ht
jzRaKstcx0H9+TU7dMo7FCuxZ1PYumcbZQxN3R9O3IZv1dFuuKMsVnq4aVhky3cOaq9pwOehuOlO
WTb6NuVAhxX2kvDOY7K+hjrUSfc7Be0bJUS/lmkn3aWIJSEjCJWrH1uz90edLIGZqVI0RgNkX04m
C6m45wupuswfiyHpudBQVbueJvqMMiHn0Vg/O45I2OiAlu4cHMGBkFrnzMggFOIgFKDq60NVBVyZ
2GFCC75Ud7S32E4GlnVCYiqEVetAtPJPPWd+DTFd+a2HXwgNA18PLNtj1mY+vWiUSvYy5DkdhwDI
VUE8Hq5U5r61M/FIno40T7u4pcBUiSyHyTyFf9vmGVbj1nYnfyViwcM8x3Id2gicBSuRWxWRlu5T
dRUHW/r0NRT6dSSUU62DGEbFRUrPv92xzjYd1pCfW3V5ENBbqz7VEsHgv3ezUuE1QnAwMHYgQsgG
aziiWl1c1USjyWwbasYLPcxbaJcNvSHyxMHDvUapw7/urP5brl3y2TeJwVLX3FVQlVuxzqS9YgMg
BGGHJnhU+6vMRkeBdQb+fKFCQXDeWTKA6S4n1C6ejVJKge4Cd5zwDGa6xDUJ3qnQKQ0kMaCAt1je
ERPM4AWSvyS5wsvoOxp97ZOOrzsk0H/iq44O0BPQn7ejvSlZ8UQ+kdCsqhX1yrF6vngmU3z1fAxW
NKqHjkXn0L4VjwF/mWeKLpUHV13qvtHVbYTQz4iVFUmnN3ufYKhbm2+QWHQHaTm3B4emDd8e3hKV
+c0GXsu/B3wxWIwiFo+OJK1yDUzCr4qv4FvdH7eOkK//GabPZqwmbrUIcOM2KN5bxxjg2VB8x8bC
FodK6Dqo0xyBAv9Ybmj2EiOrI93h3y0g0jj3CIk5EZhzZVetN9PppQLIM519M/TGDE7vvMTu44Ui
HUJr5Ub8HYtXSXdSA/qkZy5VJKHbeHlFSq2pewCbBUm4sooz0Thd7UVrO4VGNmlMj9zkgtKkxyWp
cERmS9vrLUdE/dqsHleE22TRPcLCD8CjOp+TjONCnZ08CbNt+udLM6Xr58jF8xk/EaLO1xBSXCQN
FiQWxvYII11Q7eReOCkVS12UczqnsnU3nR9gsIPnB80JKspz4QvHwoXlOyrNtDYo4QQJLanwuuXg
rS3rEm9NLPRQ1H7lEEpZ1YCHko+lOnrR/P5mQX6MkBJ9uN79dPIb2WAsdjB23+kQfmZC0ovuG8L7
43bOFZ3ivSVKXwfm00JEyU6Ear+CXOa7y64y77BBwS2MwAt5cp1NhQcfZQp5sCMWiIX5inZr2D9+
Q0GEH2n7w/udIw4+IUJlnjf9e2lxl5L1M1oZOvv44BTHlRVuAYDzcoojuQrZ5AVznOOsoYn3RWhd
Kgfa72wGgfDSU69KkVSdQJrttd1LoJLaFc5Q+4Ylr+3Yd5/FF2AUOLS6u+5/a76DdTgAdqLLQaK3
AOzMIbFHp0MfNXPQ95eNeXpU4jexPyXC8Hpk8YXGCUdKM8BubjKNlHr3y/eLJHb1NB3l5ierSQUn
y2Okn40Nue2buubeY7vZMc5GsZ1pwDCXkcE2wPzlaI7SvZo1jBooA0gNQIdjlGrGjI6h0WQbxfgp
4pnFOWX8XWtsPNPt+eJeHTF+nJX31AWluekVV82bzRktfpltrW1AkSYjwWbNMvO+L130ZIBt40Pn
eDrAyOLCeG5h0bnlQSPTvQoCVsNV5PtGLmGpvnG+NIw0VfhZcaSpIMY+GO62qQKAQt9X0loVp4ZD
HV8M2N+PVuiLrCt9uyb12BajS6ryBh0yONU7Leckotn6/Mi6fNYCUa5bkIMUhkLvMwbM5V2dhlJE
qfcxS5HD5/oYCDMGCPo19qFWKaYQ9ttG859ZqvDz6EHoltfIheQtSXOF2WFC/ALbe4dbUiTQymIi
Pd2A1KCbN45tldH7PpGgjaEnDtG2/0HIIo+S1q1o7YG96b8bi7NuvRV/P0tIm34qU4LpfFjUZerd
jP4eXnyCIw9DI58d/faegIjm8laQVMIzQoPbyablhbOw6+1BvVy0BT7HRvQAeN0mSxs/GdVWqwd3
2fiRrM2YaQrok9xDobct/wUxlyLa9nwomszFPbWNYEgNtVOzw64pR4NKmzYiYAdh5uzAa0qDMBSC
6XGyJc9x42yqM+FgApVpt/TTfp0dN/1uYi5UF2R1C6ekfQ1jt1NWjDyKHkQnXM/lDt4klLC8Vo/W
W8vSb6d4hGspiAEKxu5OMGMkwWXYlpXiGAiU16R6PpzHAuz5f52b3puFF4QWxqND4hs07drKGsf9
qJObWFjjC8GautmkHXkg3ZJUFd6oLs2RljcizKVk/X5GGRqfC8U+kcMTHujd4fZY0FeVhdkz1JAJ
QcD9A0l6c3O6Ws9V1tt0+TvrJ3cZIUcQqJrViLH88gK/wbjkgippCV1pujE6rquBySbVWRMDifeq
fPfwhrwuhW3fe9+XZ9hl6MZNSbCW8zBq3Zjv8HaQGP1q3JHt5SqzsZ0EC+OzZkT+8QQSYLTh0XJw
l6uEMsSQVAaEV1RqpWw9Yvri0H2S5t131elq5DvrTa3DxZc+9hfRkWL7OKWxgEPHf0plMmU+K0Pg
CCmGy8uSaKVMtCJWIyCuCBdyVikJkZeUXk6aDcN1mzHPWl+3ExcwlphcwZ7drQqiFm0vyobJtqUQ
nYMGEAD5b/rlcQ+Uv306B+wLdwv25L0wLpJ1pqGLRW7fqZ8u4XiM0jy8oc8aZxXQWEl/wrApgZ08
byOkA9RrHpgLlTEAlDQKwlcSsz+njaNwlOwJ0SR5v3ENcoHtdbWuLaDj8CT2kfwfP02bDo5GB/gz
L5uVaWl9YpO/xa6emWlD5L8jUtrSNJXMhTF8dNH8L980H2TY1nRxX9g52IRtKqbds/UZ6elf7myi
8vW909Q4b9CnS2ysI3uLzYlbF+tOE1bp3s0C1GLzZmdy6KSJjZzHv7Zy34BdmUN5MH7lD7MgISao
QuIudSf27MB+om5kn+BsxnuitusIMdZGj9yGKkF4oQp+nuoex6VAGAN1T9dkW1t8Ccwoi9cY62hl
NkAiEpGa3L8AWhZMF+sZZ6OX8RtluOYzudtqMKeV1RI+wswEZriIrK+FigGQbyfvrbeeht8+5/nd
DXA1ZeSPgwUkcChCfmlX/8Us4Y1Q4W+npptHj2bLj4OQTcyu6X5dhkjVK37oHwK29usoXErSuYxc
RiKgbetrYK/M+4Z89YxXX9PmsHVtkc31/TbT6C7E0WLAEj7RzZfrhrpSPk3g2icut5lW+S+hxgQn
RUPdSBr5sKV0H6LTl+e7CXDackB5VUK+Nk9Qx9FMLkBbhW1q4cYGBOb9bPDygyHNyM0DSuToVeZp
arRo58QWwdsu7d83C7S85ljyXzuxXoC+CIjD5wf9Eee5AzsJt/xFBhq0w22e7ScpQ/Yv7Cn/ZluI
/2A9pgD1qdx54xhorYFjLWc6l4fDBKs4MyW4Us2+mFMND1wpBsBMwc+46xkyc9T39hm26UBvTQrs
NGfK4rRRfiqV1YWQR181QKutbGYOJzig9np6HYsrkoR9E8SWRb+R0van2HUiis3lDHItyKg3zRR3
90ZxucNyC2fVtTY1vpTRQMryR7Wadiu2xcj81SuGRY+OB/I9OKllE6fnSl2XcL0Ma2cMbrmDAkl6
1SEMjjp7yoxIPReEJCIDN7YjUDG+1Ud2dHuMd9aB+wjNXgTzNq7HkVfX4Sa3SVl65rZNkzzZ0S+C
mboImA6gbddXf2wFNm9yF1RhOduGXczllRHu51mMmgQqzRSns+3+Jw1xD1aiVce9U5p+5nSVYZGc
J0mDue3XTEJkomRkHKMXfpXNKvHPhTf819gtXkW+cqBvVaLEqKD9wuSW2LerLCs8Ui6eJzr7Assg
lIxT9NJ265MeAnhcVHrUsnGcs/fc2MWQu37o1M4gChOtPbVNfPbrzVkzJtzcnz9zWTLGr6014nBY
qH5iAi+hLH0eDFAdDvz9H1u0oXN5H8nf4ZLy/txhYgM4G/RLB1pDveR8jIGDf655L6Xc+ZshGbWk
kBHII+ZQ3JAK19p3B5B4Z+ZwP822Qf3oLgO2LWYI7p4aQyMPTE/tgXIrxM/MDBRgxh84UJf62QoG
tN0Ct56HiR3xcehrd7xUpn+NEwX255HLoJednv/l/Y6qXc3IlUESW2frGYtvaMWuUX79zCDeYdll
8cvar2qm57Gwk64cY5R5+/c63dktqJcMx86DDYpvGEnJFSOw/rcNNJE/6M1PAy+icPijDmyYdNFy
AtBta/IqF+wPvpMkM+kfLegaVJJV3oIQKEQLAjBaOJva0Wt3QBibgmQtCrac5NuIuSNhj3oq6bs8
eKvGH/AAxCEzstA/Z3bHWxcmk5hyM9Nt4HZ9B59Prt2Fe1xWR/Je/PG7k7nWLiqE0BM+c8LgYVZW
0SP97yRQg9QmZP1CC++qGTyvN4H1cNzxAB4XMXWFiq0fKDadsOemQiuiptMZSwlKg8O7RLHWwiVi
0+IUGYXOzFesz/F80KkZTuPyEJV8inDsnnP9t4zIHNvrtEPOmnXxsXlgK38B63I+UPJpDajVXArY
Jk+Q/SnPJ268XXFeXCJFH/Py+cGPg9phHTEvv7CWeDNUqqsrQ9UezuOf+4qKjyCeB26iXaZoZ6C5
4quHXCX/ST3SuImY7T8XQbJfI1eGWQ44PCkJ95O+HwnEnnfgJNGATzesMXwIoA4ZItixtTcTd+C0
gs4p6KVf/FOoXKGm4rkEBTs8HlOWUgbHAFarYOVZ+k9uh5PqlNytJjMgNSdYY0l4UQRjWQ8dlm1T
udLog/6Bzyk2G1gGpODr1qD4t7To3zWKq8utahZnlhubasRKwRWkNzj25SfoWPu767d+hoIXHAw+
qB+rh2eRaraSkDhB74IAIvsMiFktiIBzvtX0r7mqcMGEYcTnnU0qvlhZu+oHNOhZKz1rhveB9eUZ
9dOVvdOL/iETsBenN6WmE6iEchIe9JUAY16yY2XnHifzf72oQJn9J6G1pGWH5Qwn4SL9u+1MRY3Q
WB0/ONo4am18X13t9rigpxabIFgsLc1Da4PhlWN/45Z4iediBzr6Mz94cwnzDY5fdK4WKM2kTQ95
CIb8WOueJ//HEL2v5JesNkIQK53PSVzXigasXpzrQ8ZaY4qg8S4iscrlRaodExbgn5U22tnS882q
eC0Z1Kvm8naWYWPpty/zFMUJgh5yDyib0yNcJzL6BWJSBwJ4uss3cNnv9GySZTC5BTDZPywfCEgc
CpSQ70sJo32n2FPA35i92LXK6quEALg2rh8QONdc6EA+NJnQrAapHgB9wpz9OqLB4NZeIaASDzTC
anJUDs6iWewWedwuOazrfsq1DrjcYX84XGWmaJr2/CtnwUmooAo13OhWN3fyzSX5vJS4QEvC+ti6
9w5yaiz+uvnAGg2yWMqO+vRgdCEuDLDUpHNkCEghXtTI1rHunmpb0mjBdzlMbYABspxY5wvL7lT5
W+NygFsecI+kIX7op1VLcyCNHbNuEQZvMytpb0bM/VzalYuddKSjb5bCa4PUKrLe4E5RJQgKIjo0
qnDHUy9aKYKT6wMgjBf/kFk7kWyXPpD95gXo8ew2piCwTwQl25+n0LAGLjHlwBVYW2U3hBaexSOG
yv9pmj6SRmjGDhq5GzqkXnh2ISPrDBdldBHN4iff6NtoBsiJznG+1J0vh46mJEK4waDw7utGwTfL
EOyrb5M0TXLhlOFbcvv4PtxdpuVWmZu91KCd6V7sdvAgkvvmgs/asH02Q4fzAgJMFdCFAxsUT1hL
A6xAkJdJdErIj9PdBeNDSMBdQCvs9YUjMIUBrTaFfZ4IDRYXukVrGaAbXJfsn1RQKhpOCYg/U4hF
8nwZC2x3d2S4feS8KlIpl/6R7mXD6DiAlSjhMpkA61aSS3cffKzXZoURW0WwyaQgLZkgHyNdg/ix
wYbBXOLlatVrWwawaVztR+u88h/INr03rpKORh4B9dFIVmTIfj2FXdDZMVlTd1CwLvVtB764qZsl
/gn++u9ZW2JppdwT63Tbbu96+g4gHXXwkHw9WfVqSBy/csbkPteMivoUCXE4N/dD+0w0WAi6HMNO
ruux+jyumZy9BTKhQN/dk2q/o88F8+yNVrmKasWvZEzwgiRpT4hnKxwe/UIBpGQ2/1tD3+9b30l3
k3TeyuELqzVrcXFBDs2X+3J+yPWirvd7WjxU+/i4uQSIhd6OMfAaYvMMuGaBTn7RLwOwXPZtP/Sa
U/2FKOiPi42WUdcvfMeWTQV04HnkUm5PnsjF/wIoDzY1cnZ9WxGvu9vrpGDXRMlitnSqOecEcnrw
eDQd8YzwBiT/UJGSLf6SrV5k7AAEcK8+IVsW6aETsqRG8mfAblwfVK61z4q1TkwZbdVPhk5sHHdz
tYT0iviP3v2OXbb58kvn9ICS6uCK+SrSEpZra9+IN5ZXeoVXqnYPn10KQQcEHZx1vbWIPEbrx1h/
IBG8a/s8kYaL9FmWQ0NTPrguuLpjXxYZt9SPIS2UOAsmtgSTtso2zCoYxVF688cOR/Yrw+igrT5+
V1h5l2zKaUqW7ndxS93/fYFRclAW+ylFGfebmwhXnWkfa8rieAmJmLMiBO25D+et4HI4x33uC1Yo
TdsfVy1bUd49cxwySKDPCJtw0omeYIMq40PyZjMKKeonn+I9AIpKey9vDVEyuPXDW2YYYbe46V7V
rPqTxOpeuQu8XYxK8bl+RQ5dV7UsWjyMueL9JFK6IX4jjbxyz3l/IPr/LbyTmCrxM552ledRRisM
F5x4wPcuTjEI45KwOER9OXHfJtXMrM/TuB6WHyEenAs+Kc0v+Ki2vTG0zNnULz9Bes46HblXHA9X
KycaGsI+zWKQ+B9WRhQwVyKX5KtnHy1HbCtFWLMuqnqrbY+NPgC1i4aBQCiZqHOr9CNJjHDx8byi
X03tiHyh7Xx0iE1ws3SiMwpSePux9BdRYa3TGZRZMEYuk9yhynMEGJ3XQXK/V9DYixdBEkOancvy
m9yFCB1cIm/i2qp7WfZFbJz0jk/fm09xX0mpznYpMazqCr432LFVrEfuNmNi1xpVcksoE9rMEs3r
RDjoVSj+5ShDs7oFWkLQiL4t8j9QBH7aEgoMq8mVJpt7phC+vAhvqft5ty1KyZal0IiMtTLIXu8t
h+4NnSSjRdbSw8q3Aqk/qDjw5ABiiKS0hbpditvsjmNUv0yzxL17vPJhw92Z5pQ4gwuajwuwnoL2
/hYMei00XIwb3SlsVvhSEjwqXPKKQFfWh1WBkYKi64uSXWjk8BOgJAs4sVtlgb5uXF61n8YevGID
20y6D4hsTC2tlE15J6UlzVWivHT1ZEXCpmibMnkFVm//ad5eJvBaRS6hnzAbxULQvNpJt9PWTN9M
Dz/5fOQ3nWkVjBc3F+YZoymaKsxaIPLE5aU1WXHtsmmNXollp7F4u6GeXIbJc2lLllEDd4h8DlNW
zC5eBtI2AL60SI3Tu0/I52HWibftFUBWEQjSqZio9JecN8YCawgf5IEkQ9K3Ui9At3FdBpjsIZyQ
GBxX32pd1wnNi5wR7kg8JIN1T31KoYkrYKro3+zHWd4Ea5jkGgzkQlCZbGg0b662bT8K/T/YRSsN
OmsB+VRqVvJuu6IG43v0mwvVBCzq1ABXqr2soYEmhR3m0uQCAlJHyhAwnbFcTBrEzCvoYWZbDYp1
kWutqGBH/r4ccla5VGIJJdz5X6jTKdH13sVQc64e/qMGFbztL2F7TugojDZjz48ztD17J2x6ti4b
7c6qOUAKDR1asUFDlHauhmuoerqQO18cuBq0uX/7f3i+vRdT/t6caYsCGN1btKvIQzqmYqjLHWHA
tWB0T3+qI3LJPP86HZBi/n+R+1DOw/Dk5F7cw8f6al7iE5zG5k+c0TeyZ7StzPkFqCMrmdJGrOm2
ssCX9k3ql89K7ZSDwPLkFhifH9WHGFoeWg2JMPwhKv1+2H76Engw2dt2f9SoAH36lB+cYiK+caQE
DewZrztGyfmM3SZV2xQhXg83l8qOx6MCPBPOtSQr73KLiZR4FZ/WZRQrptm7TFASDH+cwCPHUb/E
mPktNpqf3ex0grfapZRI6GH9cmVY6I4RqlnfVtngjSo1x0JhwGc+Xzy8SlT2tQUh5QHrvQXgCKaO
mv9/+d/JPtHrrMIUePuCOdvVtskCwK+N6hSrf4vjC/9NI/dUYQa2h6jr8k9/4t6m8lzyKLmUbjvZ
hh6O5iN6mCPFhb5u6sYq0DDE2R4p71BAOIoKNICFi4gyVbJgbgPp2n8BKGfH04kn3ooKoMf9NJzj
MCAxImBjlT7AqHdzLydMRSGBHWa6C6bOkYKYEVUenziCKXQqivSd9PTeEhx4vjQXyu6DQ1aEYPF4
F2yFnrpgdE4XOCVn0okwdDBTWjdgc2J8ICtZUSFhgRsZ7+kEo7Rg8xuQ/V3etyH5mQWD+v7Z0SFw
X+AW0C7bndCQPSYzTMelhjro/yh0oETDfW1PEIV9OME3UTJbuHt7P0t7ntRE3SSyWxphiWHPdQIH
nzdLohiv9VWocF4DedzpQriL0Ndo0bMMKl0OxJL6+p2NOtEyPht+ryEsd1DP0jPXU02RcH8AEFaU
dLS9afoxo24P4mAHRMcFfT3X321r//XwrjoC1aT4zVtFdrk3V0Nf9Zjl0Lln+Ovkiw8YHVX+xNk1
1yZPgzH+tzZDkuPfwKL8jJRFXa1JMzqUIJ/FKQAirQip5azPC4FmXJoIEo3IAN2W8dAJCH1+8tzB
WlaAjqAhLit7yHPat62aA/e4wiZQwxCdmTYiezvp6qVTLOncA4n5HMd1PHvqVbkERXexBVJh6VRh
JVDCcKECxVnzWSyTni3fSVBbZEV6/7vhSlUDV5lUkaqIVJRCXYnXetT5Z24wRvDtr03e9ETy8ZRz
rk6M3oamGpbv/9G6iBbCG7jHI0uJI1Q3GHolrVybYkbS5lHj+43SBEz119l1lYMZTeFR4mNuUlzH
AlvJe+/Ngihc545NT1t76331OrngxajQkKDpsd0jaqWdpmIqO2Y4QFPtEjU8tcIPMJuzC4Vh1TPF
wfS5daXl5zM3ZMBd0OABSfJzL7nDPs1VmyMjspUZusIFtvwKR9PGW4sxzk25q33t90g1vgrqNJUE
lyjCz275E5b8l50WbfAT77Q4ykYdnZPf8a6XrR9Yf0OfrBvFhf+B0gXTLjl/LB2Fr9QgR9qN/adO
XQLGQsbEqXGzbqV81fxa4xBkAi1iJxxGG9cdMakodX8eYc2jqZipCAzTk7vIxhfAWlmOcnK8MnDx
nRSAlJkXmp5vT+8s10t899DOOW00n1coyIlFPiFVjU/Kfo61AmCw0kw6GccSgucjiFmM5KW84mj9
wDLyxIr7pWR1oR6jHIf6WAqvfhMc4jHi9owxBhuSgCgpKYVOxljMLzQbZAiXuHijPITX98LoGmIZ
aPAzEdecRwaVhkTJ3FRIjQptA5UBQ1obFBwaMJaEVfXMhRPVSxRtNh7aozlsCfi4xI0g2MImGB9Q
tZiqWsuTSYl4ODgByDsX2Vb/4G4QXgEOsf7lha1stGXm6rNqZRuY/ERh9UHCH9BD6JXgj6ssf7El
Hn64mmTVYqT/9c6otqpalph9FcCd9Dt/eguiPtuAaM21ahekSGLHMc2vgCrdLWOQNV2JY3MZ5XVh
rXv03yhUm9WYW8R0azWDKcVPHyx2X/rRZWpmVkojncqFvfdtiGpSKOKfrYgszPJ9dYaFROMQlK4w
QSzsaYmXtFwr3rUIvenMWprJck8eR5baQRRBqf/SbtCaFr043ktcXaflbXGCiXRXu+cLgsUPHxAh
ZmnNU+zgfAhNfqRQNMDYMnu98ZGpg/iBjsqxmIAw1vZYjFAx/kJZRrYHielJCduXaQXL59fMlWMN
6wscYyBe2lsj/YiOqrX7DCgxCDpUX9Gp1cLYuedQztuKkzETx1v4nOEI4UugEMqa4SpxHY+GjtBZ
43DblutlEpAcIvKj93byI2EAbZgcYIE/G3bU/8uJRv8Ql3/EtWZDVWi8p8tG6fWtOg9NUXV9X3OG
fK183P6M9e19FmyIZTXWCRUMHzTDc7BeQQx2poX1H2jbHUR1d3yHmr7i1zAp7RCzi9RtHXieJshh
VQN+jk3DTAE6gM9gF4Vg7HD20TPUSWA3KSjqV00anUf2M+jHuZdgnTFL2aFZdOfRfRUPjc1dpYhA
oNtBrev0pmqYP7SLrlZ7061DcFHbVLRD9B9Xd4rhHZQv0lty6DYtTc4dNt6Nfs6rxpQE5o+hfDFa
SFr8Vp1RYMeDUyBgGivKvHvf441C5FYJT6T6ox66I2On3KGa7j46VrKXodcHmV989sb3McoAcF7y
qS4mU6wKSf2ebytjMpU+TMXc16/f1gjWDsjeU29ngSjhEKd3sbDANCKBew2HJOSOvzFkNrTWOmJj
SYPTwAX7IkhuEeFvNSrCr4oCbJWu/SDYgYHMZ6vWHn+eY7yIDsIzHohnLQWrlBUNRhQ28rg31Vfp
CitX4etgGrQsPubVyMq2EkpOhFxVbq0gNMtfsrONqSI4OhMk5viWyzGA32mutoAUVGqoQCGgYh5s
ElNmyxWIdBJZqPZwsicWiMmk4JkvLFbKWda1lDlOn3bCdb2sZCNIlrRk5PodH5sSoAKtoVGOW4GE
9Y+QFHK/7HeCtTuSQnWAr8eNzZFWWhzu9PTzwJeAX4kHZqwe1YoXfwQLSxx3ygNTIIlJlhiR389O
UtIHPcWS7mBnxC53bqsziaqjv1upLVAMhmxu7N1Gq7qJ24o7d3VtoO3Qspp5u9sLXNZR4y+5jcLA
Hyc2kJSed/xr7bkir54cZNeM7xcedL8IMHgCPtu5RKmn/Qwt9x9xndlfmFK4ypmFK12QoPeE3xki
NbHVVNx77SYbc2uTDRiJnIiNjK/QMHGqkj36O7lpNXmXnt9FyiSiahckMzTSJsPLlwdFxobas5XA
C1C54tz0G/WX5xv5alezuvXTIC3BMe1sTNB70pLLfGRLjhiYIHLJV3EE8+MVsEbuPez74087jnAU
e4NPpOKs3ozvcxzEHX9u0HAbz0JeBov3dkgubScTw78mneHPQ893swltwX11qGMslXssSCF25Nss
NQCZhXoFU+J0QSM+Omaj7rFS+VLukhV5ofIEam4lNMmJ7ZhMDKCdhm/lan+RiKmG5xqmV1ZDh2a8
0ygkn4ozTWgdrBVztM9UxtZXoQuL+rRp1nV+6B9LHrHU8n1hRepx4Sga83xt0johROVD6CzxSWDb
m6pUJgvAW6wSfKB7iMS/L5pQGQFFD4LWSpxlh+w8bj+BNQEsa4tvrSzJmUbTV5ZlrFrQ8MCZkQLv
kJ8b3arOAumKxm/T5sKLue2ShwUaKQQIruuNY/HkxPk+PwM57UQmt4evyIgHbkfsCzzUxyYU4n4u
MzIPxr47yLAlFDh0ko0GwAigXE4SfCIA3Tk0TNWNCG8zjAyJBnsiyVXUv6yreNlWOyPSOGyeqoH/
wrK1WNVwn/1KljpvgeHQUXcF+/sNIkPowKLNzyesE9D9hMjZYHzmU24fAx376jCE7CSfTNoAz9bn
C6jpq/DNv2r3yF1jLMIpniFcl14jg1KsnmOKNOvgeFuBO3p62Z7wKCY8dgEY4xK3tBiA5tqRkj8w
YKE52qyqYjU+qnF66aiMMC6lf7KMoN2aRkC1I3Mzkbkklz8eId/ZyuWHLaG6QoIqogJ9Bye58O1O
J2UBWGkAzuzb1cLA5H1aFreqEpfzSGqX/VYFCryQXHq7AxPztdKirmSsZ7sh/LLEDKk5a48eba/e
Tip4G9NNt6sDZf1FFf9x2xw26ObsNdCI5oAf9jpYWgPa/5sOXboavYMuxe03nppaYMATqR+EbTBf
i1m7cUWSWr2zYdlp6IX0H090M8xBHoFuQ5TU9DQG93FFaZ4M7OJ8bGE1TOstrhajgGuGaHAQ+jvr
kYsSlYu1+ulpRRW1bqBWJuIpCFWlc39CcLz9JOKmZDJYKfi4DQETZmkzuERK4B0hDuJxaY7bbK5W
fqzFc59TqChNpkjnXNJXn/OyeOC+BsoPoBQdQs8a2z89xusn+OfBQXoqmb6UQ36//d3bcR8TbNHt
KErfCatGxZ7z+Y4SYeRLHR+R8mGk6BxTBrJeWM7GuIOKiQqWwOnH8a3rDX0t0qm7RiFJbvifvn+z
pxb2sSc18oQwD3EPNtq46YK/k8CPVgJ5tJZZoS4qIe6VCAFOMKMlfoeGB7kaek7MqmhcTdU2UUjj
FOpwFTO0MrklYvpl+Pngwj7lSUJMJaqu6f4PNCCh3N8uk4YoVfTWD9oEhmr++Ye40o4JcvwS4sDx
QD1AybUnuybbRfyM+3ijmIAl6iO5VKoWhcqGnuinZ1QLdHc6hnpBa2Di/begRVbdWxAGQ6njFwrP
mBrda1p0QIywxOxLIDWQN2QEE7WCgXAx3lckkgnzQawclPNWZmkTMkO3e8aERyyLqFDHjaMlI4lk
FSBpnAgk64mut6+0YM7oTXtpf8wvvRE0RYQbAD1aIq/bg5HnYGgKeGz8JlBLdYHuCZOJDdwafw4Y
G9PQtTjXnevfL9yPKrp/io37Ud1Nps4P1B8uETPvROB5q0keKdhERvwG7h+GIzFAVEIaPFkxlLdf
T5qf/czyrqcn5hsJE1m9TXqW66c/KLJYLnaOr8lXbjZIoqhjpN9n7qs4XTzug9K5Bl78FTB7OP3b
MXgTGjlw2HFXbtt4SJ0MvThkkhc5mVykyKRJQZKToWw0CHhUsIfmEooZXDzImmx4m/qytZw1DsOB
yENEK06ijzOLZz6c+lPl51Ny3J71fn1n0sgzhYUoda94+PaafNoX9GVLLjfvHtfRrjrr6jzy3bul
lfxmVaPujP8vMyIrQs57A98GpRHFYeOoj7O0/dzwA6EPMJ7minHA46e3Z7fQvs6eq1CT9fPqxF8k
tJu+qFwtKkQbh573FynFpp+/4dm5yLw6okQAjtCkyQMguz7LgFjH8F2u8RgU6WjMbYYYZ1qhauyV
d08fKP4Ii4cprVWDWkbpWa4sJ9ZAfthfy3AN5vevEBK03vJ9Sh7FwBQ27hi7ypsTLQljA44sd+Mw
xhmpxl6xRc440/G/IT56g1rysBHhUevL4Tnq1sSZPUgELU7gQ5hTtqCVUbzu74yMhMM1d7wCkehr
ziPfRQU4BBThT9I9wGbOYr6Z1ODOEBqvK+T/+USM5wejVFcBL2Y2t4KpSUuk0JQE8jrR3xQTOGZz
TeVvBOMa3a+azQYuId90pvqnK78OSp4v/gnU2EeSgH7W9QQHlpWmAVdPU+yJFWGcCjFxJjP0V9kC
oZqLEjqwzgn9ehFzCTHYBV9l9StwkAOEwfD4hhKjLQuHd7I/a1W8CK3uEJh9khwovg30qu27ip5A
Ir2MI07Gbzl8GefaBEUsV3VfwOHHQye3ziKfJuH8Ci02ZP9FKyyTyWznvGPJUxIGjP2A1A+YsvAP
2ValSaPra0t3Td3bIzLgy2mnz32vtKaXEFeJsbG0ZGNJj3VxcMcosuLwzMXKQ0MuxbhrWOgxdMtC
RJ4wtJjJnl0Ttsa2XnGoTgqHC3W+imI7etEIrwi/LE3dpM/G/3ENWoVQQe52FuK+1IhWCReUrZXQ
cG1oa9QkfnEW0qOnVR4dl4zHMCJpHujYFPiRVtCHlY4a9q/In5WgRTdSt5IkVgNXYaMGjX3TmQ/j
v23JYNfpbHqhdb7ueuLlgDmDyz2pD1ozyXM5FjZyKfbooLWbQ4M9Ej5e0anwgluGHWexCHnKZjG+
KBUoiXyISiiUE6eXf3i/2oBpPbsMYQ6zgbebDIp0GgTVAyq0+trpgz4qHF4xpPVV5/vUK5DFXxIa
D3mmYfGngwXGOQgKjDpHfYE3XiIBMBw1zaGrb0WdHrg1uWG3yeHop7VYh7G6dQxU27Rqc1WLWlR/
7jkNlc6jYgxjGEwYE3+eFETPsXRDbHPPQ/RRHPxpumq6S6S3fqjUhGIYh+N+K0lEcT68jMjXdGOr
6ZFLfUhIui/kJopKrpXQ9YL3wZtZQNllbTYauniaS1scJG/Sb2JSLYlieCestFBLaxZvRpSE2XTR
mBxFkARhs+Pxr99gdLRYT1ED/mKVzT80pvveM8TtudRn80/Y/DTrxmITWpvmp9hXkTZx7kK/vMJI
j4IbfA3FFsuXWfAnOBaLr1FX9s+6bcUZAZi0HQ/RP9w1xbLF6ZhsWVZHmN2LjwN8zRWVacayeaGb
UVYXify9498LcIp/oRV4IBb3XIFQiPmdnzhqsvDKJjxqvdohM61Tu3o1midxQlnH8hnCa/CigU4t
Go02UHeFxkjqVcanavRcV+O60lvBEXsXUu9vZ4wEJ5Jmj4dvzyPkAy96+PI1VUixS2LcWErrKHGo
pQd1itajU48LtnDXTVXB20tQ+krz3S87I0n6GSusjz2BlxroOPcI79hJj9BcIhQLicIKBxs+ZVRl
Pvzo2dFErDT3HF+sVIdgnA5YOrbDtSHG7+H2ovHxd2exyPkX+pWEDrxZHjJf9Ju8ubxb5h1/7q+w
x+SdPiLJCrk4Y4kWoZKPxdP4ocylWdrvw93ypXlf2ncRaFz2d9G2fW8B4DIa1P7wABqfmem2yksq
bDYKbjgd+/iPvi2unjc0/w5y+MI1gtDiiFe0JUcpgi+W/qaLxr3sHPAKGkK9NBrxrKYwpHKODybf
cqAhAytrjB1b2duJExxZpnoXlUgDEhOay6dTBsbZhHSJ34u5LKYJzGe/PM8/VEnH4vVM1Yfo73tS
yi1C6OZriJMX2PRv+IeDW6ih3+YQ6HPulfHBK8CLmYSb9ZWqmge3UWR20s8Sn+Fkum+pphJreRoV
iIVPf7trjxVt5JrsGSkZXCBvAXXNfbcuWRv9EfrK3BJcoW7v/+8IxGxxUgFBENatdyjez6QzDGIj
uWXt2g5J8NzRKtr0axbIho/mcFOdqPSCZuVDLfXNrO5HajUqZD0cP7WfIE5DPsgV+7Xj9wT5WZLv
Dhsh4TfgGPR9JWUjIeYXWm8KB/n9srBuKbBsz1d20lM1iADWkGGOi3xapmi33mkL1LHOlayqRSBr
xP2rU30fZRi8Es1mYHdMxUngJKOCe9tzmDQtnK1oknoU6UmoMn587+7Lz4cTJNTqyTr6JSV9n5+b
WdVztObidGnTm1qCJ0cgmfKJuPUJX9Z8KnUw17vpRJ/Iv3zJk5gt4HnvCfTl44se9lPVRnF3j2CU
bv+JTO182EI9SfIIq+U+m6kKJLMVb9348bMHFSq+b3XPTanaG5nXjoWdX60mahzewMdHKt/XbvZu
v5IxZjvW/4eiN8aCXQcbyUDqpJdOT3DR5vXQtUxKO+ZvuqHUypYc8aKefctCg5809T3ELAvw7asT
ADDIJ2X3DylW9U3bbFI140IwwWzApd5jhFynzyAHJt0FfXldt8n7hcFr5VqEUVwz+07wW4XBol1f
/XAbwQnnzkY/ZGIGZdMEJYEHiiCbLX//BTwm6gmWjcUFdraMk8oV93TuIjL+5wuUUbkD1zHhzSRu
5hXR1d/sGZgRIZdFl+7/y2+g70AZ97DgNX9XevmbUyN0mi1yQi55wdJoL2HrCit2Yz9J5PhO3jU2
1Wq5azBnYI2t6Neh0Om1ZJeuWmLgDIFb+jzO/jfOitBL/kLImlLgCE0KfBdKoziuEbwqsZ2ttmuT
aU+nLcsola818SFyds5QupZl/ySnOuGmvaiXm9ujywPUR45o5JPPeAamuHjwXYBNZNrBwAXnCT5y
1VQvXyxVY7YMutLzrpuB1ygtNPNbFhkPJI1Q2dcVU3VYNnqwyecm9X0O4ijrtNJLdWlKs4BD0Gyy
VhsizTwJ4WOw1e6kV/U0bbg0QZpAA6CNkwElmnOOYoT/1kETVstDHpXm4t1IloKFSkwfkiDO/D9M
QbwbU8wvHmNQW0icKQRG52pRS+8NUG3pvQlHEzWBIFKa6S3iXqE9Y/nb3tw5tF0J74BMV9ihrWoR
ou4IKTJjLiaKfQFmhCtqZ988DZcRgV2KaxINJcaOwkIP74iaQ7abJAiuECjXzZ48s2ln2pKh4MMc
IID9h99eQAm5OEAEYbcaCVpBmL3AUc+VkfQa/vS/IY8sYPz60uZ7gOc3lSj4GZm1EKxV6vXDi+zv
cdwfB8cCLkCnWevawpPk3KhtZz5LiZDCEojy2Eo8HAtV/SnddxqOa4QD8sSkkl3/7saRXrJsXw6+
0eKLelirZPpC+JqOBJo+E8kKkH+cuC5CjTG3+NM/25Bxz4Lo7m+hP0NRgh3LwIJh5FARCi0YokJx
d4C5LRuFgTaRR0kFODFbUaGX9xXGtwscShhQh5OLSX2U4947yhwEEjlqoDpj0SlaNB7q/Qlr3XQN
SwV14ukEW65ZmN1kb2zfvJBhdPzmLEWNBEd1puhl5A0z8CHZhiPFie7M+hVHqTOeCmRaKDj+FTS1
fRIHvD4gRZjvdAIMjnO1IhF6Zs52QmAP8O9ROrS/wYEtyXyK6jLUcf8wTCAFkJ+wCt+Y9DrslaII
brw9LLW1edwUhBIiPoTDLB+pwj1L7zNEkDc5TE+a0Ldvr7o+C/dQgT1f9QaT6diaxB+cio9ueWq8
q5oZUYktO71v42G8Kv2yhrT7gvoaluemODMpNWOXwKQYk3Aok+FLyLLgpjsciDnm2uTdCtlj/XzD
t4+jPZxQfq4Y45lSJwnu4Z17o/zwzch0Tl/CinKkPX3O0Rugbc25kFlPJeJbbYZlXmdWY4tQIpCH
N/NyXK2QuqlLuMbVZpdhKB6HOdU+MFTTm6TdUY8UFyvYfuiS4Sun5SM8QA4HAUlsw1wn5XEbVXlx
PaQjlhk0JINznnCFyfdT+FnrlVLsksi1gEobKmTvqyIgihNeBgJ9LXgRKVv/ylu4PF4sGnqskj35
7BSVFD0ay+iTHaSCi2o4z3ieTs6Im6gdmR5QIdpgxVwYJbxoMNZE57dYvGIccqkXuaZjXAXTqymL
81ae4oLSQLGWuhkMn/fkKBX84Sm0WoS9jFJw+iFo4FBs9sIAg/nPxId4kUVEwVwa27S9g31xbJld
7NhzkPr6oM+aPArgTZ7zYni6erPS+h+b3AXnDeTY0U+5ddx/SnzPUqBKHixhBy6CKspuzkarkdCw
jEnNU0VgrKPvZ3F+j/C6iEAqJ0fuIUj+3YunX4BXMLjRY3/Tzwf4HuNJfK0/Zoc6uFOdU4gkreJu
F6V7DhG+bHGqefx17Gym55iTGn16O+q7u2DlYbvEgC+QQgYLOW+c0WO/20STOz5xps9Y4jsJgKO5
KAT1TGkjhFFY+zsUzy7xIQ83J0pRX9MJ6GYpkYrpwUkEpaoqsJAe5Ix2R7IVpFXhWnDXZ5tuervl
DO4+NFVdk7w6vqdozfkn+6KCtGorM02wbXBgXTYnzhZ5c+qkKUv9XVicDtbuR/WXkVRq+PSwgRut
aR18SVjamrRCACi5H+ZaXHkS/jubVT5Z7jG/diciRg6doKlvXZ17kmWVGGxRkZ9Cj6V0vbc35JJ4
IilQdmp02jeoOCETwtIZyjB+6HggZgXC4IlC70cEMpJUbzZpb7hba71XH19wd+FQHfc3muS+ufOG
D3EIveLZRDGjjxJCxvp72ANzSzA0HTgswFGcdXbKrZr9D0RU8K8j4q0gZqkyI6dvGeKoUVNpB+Ia
UY5tilUYvEsrYWnw0ewCWDAjfQlz6ae2zwNNbk/Ysnh5Z1PLI1t3vaNGnJsGV1f8yUAH/Y7yrEnC
Uk92SunV8Q3TLxGllNlAbkZyIkPuFZtLGxErBHf0lEEtaLzpY+qKFm5XGGvxlBu+P/dhxvE12Yac
gKCXVOJoUNkkvgx5v0vUBxFUp22FcFYQqYIAfOgS6N542XcwEMxF62K2uJ6xjJcCAPb7t8XLyrgx
I3B24DTmG02tyHo08oCEilBoWecjDmqo3tYqLlplyBJSvS4KR9hLioAgN7ojCJHxgnLYJm4tx2od
Qdq8blYDU94UlmDYVfI/6zjkrn3y8WWsZQc0QQb40PCuuU8Ju/heIzXSL8blZMoYTFpA7wOlgaP1
2f0IVs3S3ejdbvei9IUSE2sd/Woy8xZNIy4HcX+h1LcEn8IHfiyHfYT4/S0+WoItbeh1qyzvL+SS
uHRm3dLb6yQhVoDWYG9qgbpWV7RKPmIfHyfedzeU1uS2PIwk+MeDV4TLWL1I/irG455SaLl7WDLB
KWlu101DpPItlq7BcIN2pKqe+JXBDS8UkhA4Wuips1t2HSzQiCB83inF6aaNrN3cqROvP7vSjWcy
9SDght4Gnxrp8i/S3HWM5I6vLjfPON9Ln7LaLBMhbN9T6KxFyXyRvmgD7m3BqUiDv/z8GlkboS+W
0cnUByplDWhCfyCV//4if95S79cGTvfo3y7DuKO7q9i7KfIC0hYukkolQr1+12oYSn8NbaeiUK5p
Z0OhyTWXJiTHQ2DmmaFWxeAzFEjjlbtuWI6W4CYnGEtl1fBCGvU3dS5oV/BPBQyZZPxmmV48Q2vK
BFHolpabQ2yvWP0wcYQwwx6zksk8G/Bkt6z26TNtB7SKCtn+vAo/wRVDPCinWO2DUi50u/BpTA9s
pkHeDnhtel6T6dyRRlYJuf/Iwylf04UzpljmntX7xGw1g0xEJDy85dl759yvNbDtMvSXuXyZkmBq
zJGmyBW9wDKzPMSI317JOnZ5TI11GHaVMPsS5oOfht/FvvEu1nSk5VvGCcuPXmLE44g6vvCaLVyv
Knn6WivOCYgcU95mJUsRcgoIiNto0m0q8Y7BA5RQJzkI8/vNyLX6tit0fLxsjnjas1xa3JWj7tXS
AW7osGVcmF3JSN1iUzXW4lJh/R20i/cKU4xCpvfxbmQ039znI5vzzCQtaSItUOfXVvHMs3bSOFse
ar6x/718o/Kzz1Xd39nbXKRuOfwoh+Hw0OZlsy+Nu46JMoH5U/XUh/cnMnaPxm+OuXc2+i5OE77B
CoHbJAwQgogxEzxbrcNy6VPwIGvkXigDuwt3UwkNJC6Fmgjazn/e9Lmt511PgiSmlsSQJJ2KWABa
DIiqNXQIfi/jMT+a64cYB9Q9Ac24+CV86UQmmeXDJ87vYfk4ZFBe7CfrDbbxBcm1mZQtYmU42B9M
u1tgp5m/f8UjO9wYOZakIXKMOZz6HIq+QdC2DbIQg4bWu7BbhY2al/iLH7qs4/7/yDNWmiQPztGS
qTCP/PschcCcaSvIbrHJbIrrn9ea+qm1pQu9ovjGZuYWQseg7dqspYrN+G5dJGqN9pGLVy/aM2Fg
YXawrVzIK4kZCPezmZy2if2Uvq66EYDyJOC50uv4KVQn6ds4nD4tkj3J3SJez4z6H1IAHRzyuMu1
Ipb8UjnpEOzdy/qSYI1Up1kZ592KQOvqPKGzkCTiasaCKXM5A74C87LcQrENhnDDE1ukEezuf0GM
Kn2Qq3Ol/CnvIuhC/LLfNg95LXkw+zCED8LtdqjUyJJsnwW1gIBnmwrHB7ZOkA/KXRwjLOdl61CM
IkZ8wvc92dyFw3UmhQuiZq05ix+p81YdWndycM/kV7FLU/pa4Py0/xmA6Y008AHnAja64vNTqYQ/
k2kX3TLyfdtrtmYaJC3eCtxY78q3cSxmuPgsAgxj5Z7EbvWrNX+jvyJywEQQBU0tTWFQCUE4rKMe
G1egQCmN5N7nv1a+gTHOn+5P9KUpA22oFWd/IyacTbBhoS82Vvu8ow2mMRLSywUrzby7I7RFZmAF
xUhshcyqZpvv/i9F461+lZ5uhbwrAH3ToSppn28o5nYFLxaG6M06KqLfv5GujZFekbGMhaTKrfUt
pOunRhX7ZXSI4V47Dbrykk77l5TIUOdpL5F7HLDth9wPs/k8itjHW6YTVmlJNnE4pxuvbkXHaACt
IR3IHpYnvgAksGK2ZNwvsdWDXJ0/dmhuvhlvFRRyqC+CPJCi9siUnk9gT9dRo+mjtwQadKkbAJJG
GZWN8xcZHuIYIAyTF0NJodhyJ0kSA50wkzfLC7+8JiG9SOMShVmQYD6ndYm6/3GYRwPLFnG7dFOy
KZKJrazrk4+7oi6O50Ek9kioSTG+dy4R9zUislz2EzkSrXJbHgeJsw9DphENqHXK6w9NcqIN3NOI
NDCSGJ8sGITGjtQjaD2S5R4Prn96FRcAvRPFe1wLenI/KJ37vgShqZjoPxEQmR4kCEdEhkrvwI6M
zC1Zk6kyaF1l6Gh+IxQF1C9Oo5QFDNiKqmHHZlhk9D5RqFMJ2u/SBIHwD6ZVG3fFOqJR7XZ51hxm
xQzqJ0epsZJQyZQWAQFAXoJxbPgpg8LqTdBgguR0hojbTlOwR20byDo8y2JGirXp3wMq+b6Jw+Zz
HNPy2napO5nL8GfhgaWfnrsZPVVky/WzH0e45EnEo8XB7pQ2qtfo5vwP7ypi6AIV0XcHnhjrjr+g
VlFE3/HhU7H9p88C5vm6yPHJfkUq5KHU2gPBSPs8zblkri7Ez8qX0mIWoeUECHZeaKOUPjd/Ww2T
3hVE6V+PxAo8m9wm0cKau9j9nOpFrvt+EIRNkBatvO6eIrCBWhPhEAheU0xT0BNSCZ7VKQ65sXqz
r50TYQXPFfNOq3Ya1I/0O6NljNJmT4fX4+Q0Gn+5bJeHq11MAzI3Zyqi8KSRjKqp9dIb/251u6jH
/SPv+ZX3kDn4Y69UjRz64Nrxx+kU3wkjGHXQI0lmXG1CkPn6wmyAc1Zqr521oq7CetyIQRRPSDt0
qrUEdAl9duF6UndugdvMDZ+ytJF29EQbgReYmZEcZFerfRmoArZB5avH9iD1CI1zh9mY0OnGTafa
UUx7dyAIdJ/zjNoeQNuX3PKEyrXrJPvDZ+OuDhwPOAcITeB9/tmLulzwgMs5qTWpPE0ob+Ger13+
dr2RmD14VlF+KW2pebFYFgmYULMfZMDRM40R4cOSbWiAdc/nO4wR0uPBqYkEtYrVIE63mf1LyJz5
QLtHY06VzQtkGUGCfaPGeOInIm3W85OlxV9m8GoNOWkswqw8uFhze8uVUkdp+v0ctAXLSBRzAFpV
qUS4CphoMeeI1aZsQF3rJaQ/rlfMzx3+a6YNAvU4KDI4sk37xqkPAm9OYdoVKGTLg0uWJFQFBIss
W8TupCmMQLg2TVQKSPmrVxiLHsZkTEKlX5VyCA2+8lvuFm5pPauWuFTYE7Ynjh+fWxT/Ved01rj1
vu+zT9/bBf2fagiZ1lcjWYkysjbUQycS2XQMq61Z7d+h5HBWIIVmJlloeQzdFuM9HGwbqeC+0GXU
b2kAefYm4nX3FXNS78JXavWnAjuMpWYoPjRd+z1r4Ai75aA/DzwVErNsbqnDAkfkX/ffDKj69dTZ
wAwPKQxzuaN1rVUHv6OCYFK3vQMZ9uJhKfQfpxW+2PcmslWe359XXsUjUIk4cxWdLorXja4qumc/
K4cga7D642gDGFP+OK5XiB63A5Blm0Oxg/7O0FYzO1f5pUSCZRWDiueqX7Ds8TL/rEaGzBQvmB2x
DjeMhATIS12Qfs4YDwi9K2NrbFC8DyQFjFlTYxzwyQCiY2xmbeOcEMc69GzPcpwY1I8D0HeFemAz
pK9J6Ebk1d4CcCKHo+ynXkeflnv4VOSZNawB9DZ3PrElOWt13MslQ3ifNKENOFOPacJcLzlZIOrL
0ZqVqNPoSg4D1zBVLeDufE4SHR2JfwqfeE6LmQgs939Lcdgsv52i3lSpLliHVEs7CU09N2duUIeS
O0635UKXyxSQt1/ltp0VEy2C5RihFAHctA+z3p1/Zb0+I1q2eanWH3XYBu9souWcL43oUgFsMQo2
ixBw6JHv42Mm4DND4X0qMn4KIMn42JBLpUjDh+nUJohnYIDBSBiiMqcTAgnd5hajK91gFL8JZZEV
3BBcy4cycV0tau+GZhioDZbfO/9VBSmrgMZYwPSLrm8Ipp/MgUcEQxwGwsrxSWACWOA++LtdrSDu
zl063xNFrjJ4iXIQw0R8gVWu0U+tZyXYtCswU9GNMYIE+R7jRsQY5bDyKfrWlM6WgyUEtjqRwU64
uZtZlg+duIXygcAO8rw1orLXRM1j7ZV7BsBCdOSBlXr1FQt2N8x2zVFM/2R98ud84RLXMp/6rcrK
JR7ofUo+JovaFPEVQ0UBpNC5zRoMQU6RPwm+qE9BmrJRRtWxkNaAwzilarFzUD8HtZUq9pleYXaQ
P2SjAAVlMHbWIq7BlSxPultjgPXFZH7Gg4TZgwj3KULagISxUVXI4QIT0mUiM4tlD0ay6eFFIZrX
k4TGzbVyjHHgJD6lL+S8w1tZ3GggoQNVpI8/2ZKMHei+2f2vTGK7Cx1RMRkH3L5LCHdF9NUgparN
wxxXgFwOak7DzuAcYTrAGQRinbxtEPA+A+atQswusF/Sr1l/r34QIYcxAqB6SqUrAD9Osltpe56K
pn3fvKmXaeK1LNxo5xYsEgU97n/z42ju8iWd/mSVNbhsHS/p2mbU21Q/qtjRF43KJ80ymiaySdaH
tza8RamSUV1zv+5cxFlHznB00u3gATuoxnh5zcjjEU9Kt0+iZJDV/RzMcAUxoimDl7Qimj03b2Ni
dfkZ95FkQiiiwnFtSPoSXUzlSjQGc/Rpajg+Utf6Sn0jRsmSDlkpw++fzdtf9fVk0h2Q2tcnNUon
q4lW/VnGjQWNV9z929nT/wkSTWQMTEfdrQOZl5/rK1buDTkbJ+QdyYpYnG8TMUkQuldqLcIMcU1z
upC7K6sb7Tooq77ljkqbVf/yapv/h4e443KKkzyz5xS2HjpRi/Woi80ulpAyyCyhSJpYWous8/8j
NzYr7v9U2NgmNCxBsR18W4ALTZ572U3COzN44BLSwN3vujKGXoqfMvKWx+xHi/dzZzH9IfYCOO0j
FByle3/0qs3lmzOaqfk/8IzjmDFFo+CfRE4vsiDQOWHqF0rGbA+nraqwcKCL4aSB+w0QNymwMDB/
ojS5xq1FrBucXwPECWf1fLnwEQagtx2c/nVzKMJYqMaZXWPbU6HI7G3WQ2VN32PmQ14YNlJH+Fm7
NiEIVirM61Y8gEo+kabUxkb/3s3YNd3Gwp+XUHWo9uCu5PfNKDrpyrc42ZepgXaC2qsfYTitiVP9
urpLzUH6mT4wCS1dmlHNZX0/QKF7aRyRy56ODV9hsh6Lwqnqk5k7ANTtbXQd2NUBydCesCrcZQgA
DToGpeEDRQHVl+iDNPEp5kB5AzS/Kl3LwJ8iSSBFSyF/CURVnLEypMULjzc7NYAmhh2SbmvqnCzX
XL+E4X2UKbevaqNP1mFAR3j+L/95NQJGX+9uvEogv8uTjXaVazWV/nHMB+MJ/3O+TgM25HtiTkWg
AhPvyKsIHoqTza39g3j7WUzElCJLHIe4QrAZzzei5doX4h7U9/KNUaRPh0od1/17ohvabevRjJJB
kgstJAY5kSiZMmpG+qgosjf5bNELB9B3fraXOXz4o+IsCQGe+CEnrzaxwAhRgW5Nz/Sfftvk/6Ob
cXsJkLnUT93maiqpLpeBaPQ5nuBwU920lfeFk/7v7Gf0MIgQSlVbwthzrUkMugUC3h7w3yR2PmGE
spVE76qOutUxsxTWiTnWCqxKYjWamBw5BWRdGtwKG5k4Oha9WyPy4paQcj1C57IHxi3yaaNL+UbR
gxsMS80W28Gq2Phj1zLWgUX4oKrdxf0A0XGP4CvsE2T46hEfr7WncaAS3r4LRYZGtDIwpmND6p7b
fl0gE87hXwOvJX3UuDfpCKNcembXwcpmxV9qI8XW6PD7wI0qilMxUtPZriFnud45oW3JDK+emTD1
pxV4OpTsBO9Nz2BnsjKA60bYs0fzkAOaYfBqFFW/vM/twWRnx2sGHyXqrMP+n5lAvFKPUdyNSmhy
KcRHtWit/5DhyNyL79i0elkWzqbZ54RMaRf0UiFsrnCpjQ0zagR8wNr65X5aN8lXg5MWH2YB7fjc
8Fsj6a9k/2wc4m7l4TizHPRiyrEV4MiWX0Ka9+kfHylx5HCwMHkuloVV/xkpRtqzPZ8mBtLfybiy
SrbNOb2w5IPNkEjIcIFFh6bbP43/BAFg7HPToqLqfCYwr202Z89C86ZGppJ5xCy9zwp3eF1dgvBz
xBQeHfEnIRs4JpTdbISrVK+VI8X301sgDwxD7hYn0sDUiJXMBHyuGnqAUg/VJAzcnxCO/+wyfAYn
+yiDAPeNzkW40gQwuZBb9shrAdNCv+v3jxvVpSbftIb92yNzQ8At1N41SnXI0ryAYTyfpZXZguh8
V1tVdz5LZ3zoFG57FngDBNzJb1oMPhiQwwXXLcyHKv02pVzbDh4Eja9EjAeeTTK0oTNsJnKjcTCI
6rY04sd8iMzcoBs4Fq4SQiqXiwDfECDEi4Mn0oZVyodSNbLb2thpCX0nBjOA9ditROiv7ac8U5Kj
eybOv9Nvo723/ZI2MswNxuxMO5fGSyF7FM2qd7cVLlc1fdm/Wx8u8wtvkKKjsA18B1bWTr1lYBzH
Avg30953K3JsCrtLKfX2uQoDx8rcNRjdAK3cr1SKioeVNhOCpPkKE80j9wuD9L0nSRPeWNO4N5FD
TN4KxgeALxPxpNb5Xcq7jEgs/0ocgpkVzyvVBdQBhZaZukJtC2KVOWmJtYSWBquXB/tSNRE9KaRC
W8AIU2W6+y2NraLY1YWI32SckBAgkiWOywr99VttWIjWAW+6UwFtm2Rs98KGCWi1yPbwqVkNKzoV
Vy+K1KfX8s8Xg7pmvXHNL8fkEFWC+1I36lrKZTtMPPUv6beS6LPTa+NMRkRrPKLJkZFaLQJg2Cea
ZXJ0PhNwMRqlOSOL0rrHDSvVLgiIg7+vfpUGKRptN5OMc7U9tfGNqTrk17uaugY6hLA39MxnMk6Z
CjUDsKUI6sUFLXCmzA4N1GMa/M85VcjvZADwkzrSm78MlZwnABerYgEigtWfAaPd+jW3g3JNTTSM
TYq68iOvGWD83C17Kw9r/KZ94XMRAtsrWEmTBc/qhWgb6U4xH6TbzFnVsIeDk/9LQSTqkGZXAX82
rlSQ6hQa/cBB7F1OMgKdQW71RBMPCIeUdiNW6VHZg5325GY7GbsBR2dZ3mL+Ec6aYAZBtQAxzt8a
n/gImbzBRVgzwUb1bx5zehLlu4J+xCAA/UmoAYrXkiVTKcn/2u0ZWSdc1g6LeLa0Z4DAk4/nCS2v
sF27I1EjhXalVRdV5KXfG+hjkB9kk/8MjUJQIxrfv1E7eHytzus1mtgYhPyw0yJjbMALK9WG3tDo
AvEZ7WP4BZN6Ul9W/xKPB6kVR5eh9VgNJYuZsXx80KlcJbzhWybeRiR3CwhJS+Jf0q2l3P7Lnh1J
tGmaLWZMseTB8XxLf5NQ19zFrmMfBJ+t7SM2SpACAHtgAEEYG8rgFP/AETTvpjirOe6hFhSRomaS
T7nVy+JafnbA+dFsE4sMmP9x/dSkQVdlpRhQ2qCPI+W1jKQpt+JoDjUW8Y+67RSV2Jv2SLFjUEOj
1fTQe/Ey/EHbkSDIe5/iXjE/vSSun9LR4GT7tcjlVxTFW/FKky9jCr7J/bEOpH0KMQh5aZlVo6nF
hXH6kHHHid2EXyu0rTXgO1ASkQXzypmKr5KvhPqL6cTob5sK4WsQBhTqj8c3KOJAO8Zc8ZwT2Y0z
xtRHKoySE0O1AOm/9dtUEl1zZZ8Q7CQoLCthe4FzwQe26ltxXXyv12zRD6MCBZmh7vOHryKmgpsV
sKb7/mzx+rlmks8OaofQsuaKm0GBgFiu+U4wJZHJlClWUy7F+UNtBFML005qTTM6RNxpju+Ef4m7
diRrsB4hNLhkSpIPT00tIgfOulHF7nlae/Y+S6QX0fCtjlozMESLpz8itXxW/xYUbPXL5TVUPRMB
BUTB8LERAxvFO8QOFw+5x49SlOCmQY+14brJM0Upv9NijV+6vqq5KckgHRFv3IxFmEAXuyD2mgIc
2dx5P8D+I21xzBH5BortZK4LN2VAhYRdzJ7tjZu4fiQWMHvefJwCHH+ow79rMHaG1dTSkjezSsIz
097brrUp4BUmJ6XhlA8y74fxpCkT4izxt7cFq4vPQaZfjQv3zoJNxj6aY2B3oTwoxND3nVZqcAww
GMa1RUJ4L/6GM/Kb9s7vTm7daH90SelK78dLYIYIeg6TqEFEjx6mweab2ONYLtfcaHP7bKywU5wC
cBrlBqF99/ObcTvVaTj17IlMrcHqRZeJ4UgtwS5wmQt4x2xPKlY+H3BMBK2aAJgcm8dNZi/cNkMg
45NP97sn9mVewuLqL+cFh13SXodf3BcJH0cAVSwciyUU74pzKgIIqHqyjEQn9oOYpwxWvylr7dui
/XVcSEnDVW/X91syhGZHH0CWu+FlO0U7jE7BAGy6AXLTzDQ0dAYtRjgW+dKNpfpna+nY5WRtce+A
PmhqU+Ts+VAtNRFYlhvABO6uqXBZnZ6tll7iBlSB2COM6rdU1Lu+o6LQBtZlOwvhcKeiqYtL1r9a
jUGwuYUPcOvygbI5hltH6krRahKe35jSUVxk3CVs7MX0BGIv93hQ+YJm4y/L6B4rKsI5D9B87YgX
Q5opY8QNzLowtcbvIXiTvH+Y+LkHxNk/2EU39ffaDiLF8o5TMnMWZtsvBwyOmfYcNQWR8xUjVMM9
Pg6au4cjaOSf3qY/iSn7wIyvj2Kdp5zkCUiNEfmm4GzgNzl05OLPoFVW2gODhGgDciNkcX+AeYT/
XmfKrOSyFl7nRtB3hIb82RcvOdv8+JdX7L1arBPYI+0qvvrxnx4enGwApTqHZmKJXfuijLKRp7A6
HcUdktCrHHYS4WFUTTrQ/u9iRJhjLsQ63zAvbL9zoRDHl0xvvTy/sgiGvSIWko5IO9UUQQ7vKyVD
ZweDVa/Z2DUFFGCGWRTejRy44HUombDjMJgfTZpB/YoT6m7MNB23wO3DzLLk+lWC9rfmpguZd8pm
/9uNSCP1zSPkROFfa9/JcQpJ1cnHnAxG8Cd1YuS4kRNzd5xQIF3OwSY2eOya+lrPy5b/Z2AgP20L
Vi21eGVrDDtD2XrZWI0xSyy3KUOBQjppgtOVsjYqB6voAhko49c5X8eUHyrf0KPO2E8XLjJsFcYn
YOMrTDkQPhmte14c0dsFczcXtsED2DuQiPNmypyDBjEujxrer6GXE1svzl4ewPXrl0imfaGx95GT
zjPK2HXUIZkBoSitaHiq10jDk3Hr3WWmfeUAXHLfyglqugZzGoSgEzqDK2S/RbdQ/TXJt9zITvae
UPYzC9Gs5wIu9p+4VOZfxu7Djos9DDfDQk1Z4Jg95uJP1TWPPHnYgSaXzhRxS2i7VoptJUpjOsf+
JM6XYG6GExb/t6Fs2Dd1Va0bmTE7sAEqhFgdvSeHGPHiyTWcvyMVZ7trdRxlX2i0Nbi7+pj0TaGU
Fm/E4l3ireL4+wqwekfXLzBUYdQkB1lRH3360r2dpz0XAHoLGOAiBGYBhTY5HqIGlShE4TYiyvG2
PzZCezhwuhrMXngj4rz7nbN+ZBRNwtPAzohXRLjQ4otdQ5f8mYPo3K5NwbvoBW8UP1HAnNm1ppEB
InEdS8rZwOirhRgZChbaqEngtNNGwZ6/aoZ2/OCUtLoSF/YITMRWERNLk8VWiTwMICDmxiCg00gT
iYQ+BWvcbtGxa3H5MXO0nafB20akXZxW/aofRQhT7mIT8HMGQXBUcowq7Dr1NWsXMKUEJYZ7bqbS
oRp10Q9Rs/nU6ywZksK5f4pJjTzP1m3YE+wR1dDiKPknoc2L8z8hF7zvfS+BSGv8aScrbkQlNSNy
Jidv8Rp+f1uhJ9dcKlfiZJIhKkuXgt6xYy9xD863QHy0ft1b5ROiMZffISeDYGcjMGlC1ZxEnYtd
P2r1XcgJDpT1dcwVbNZDVjY+6h5fbQzEG6C+RvuwjkvfMtM1NoRH/+4ac2zGPAWyVOp+wIlypezm
NUQqWxZlq6wjjjuzXyFFQ11n2j68+3fTnNS1VEs9tnr/l6t2GPC9jsx2WMyA2tTPnvVWR7FQ5mR/
pRZJNE87q9K/tNijuHTuaRexqxHu7g2LP9a6TPI59a8iqrbS7QuGFIIbeWCvYurjFKdlvLv3++Xu
4e7xtjObDNrumeSkHxHJMRcoNGqC//qDe6w7XrPp5Pwj/xrd9sii0vBrax5sPzxDPV8Tf3OYBB6p
456+3gn+CwSGHnmq2AOE6p+YmkoTuu5Zab8lq4Td+GdEPTNYTX8QDeRAJ9vCvqlegWfoEI8SAYpS
8/IIQoFvrFjcg1dcxDx8phXd9kxHaIx+cGoTkU+/d82FHsq7unV1SM1KyireZ9jjTqi3/ZAdo+8I
dK6hKUST+IlKRjz5GMZizak/oFh1ZtLgYS3zl64ua54PQQnNhvj5ZFbXKHCwwO1Bwdorwh/fTVxb
v5DsGruTA4pERu40UOWc08g6K7HZj4BRJXmp70LuLOVfLqXRkhZK8v5ebnwJjgwZgtqaCgbiUR1x
VTVHMslIsMpmnxK5guikRwsDdPPMQUDot13d2Cdqimnr/QUqI/K2DidwrHVdufaaRql2zk6FAaHc
UpQRkXSexfAGlU9cb6Zkr8l3nf26AwBls7AFza/xa7PHC+QPPhuF1pdAt/v0R+BzwZ+pCxt/4NBE
sGhTgpLHmJbc/vCXvGPcNCn/altJxIwww5eS21fXRPkf39qsYRWUg4PfkHTc/dcWgV9BbewLfDTd
ZHbBKAl161PCGHZkGOPPZjmHyrjus/JJy4aUAkKoF5e2lHN+1hFvv50mVU+PUuSohj8lVYRdFdte
X2Z921IHH2lWXWm5uzi8bhXlwG/XR3M/feWC+ziM5nVpWTwOSDbdjKoZSXAtMWiw50vrr4e60mln
N10FQKtM6AHhu0Q4Hw6oj50mQ4TdFX4mvF52VjVKbh+ZEXbHWozWqcWMuJcvOVrN/sKRT0C0cBIe
fy3C8cnbRLRkTL+SjdrmqI/z0XwF1LXR3h/xF04MKmVxY+IwrhSgNzBD2ehvng8/9rEM/bmTaWe7
k2uuiySr8SYvWi3hdwxEbg4bML+qrBGTvwg+SdSyustEBxILSVtZiNuTmu2c2x7sXFyz833WAmHj
ls1DEiBoGlGQK22QXMrt7DblR3y6kuSTNVa3i1F3uBbe7b/lLLPtw/2zyc2+YNhDcN3ieWZoEf3Z
QM/7zceNZuYkS/Xh8GM7ksEfr8fkvv+l05F+sfNhWEe9y85ZdDgOgv2REOdiH+4TxiB7UZxKZEXC
yCDfJnI/NVe8rt9yTxjpsXqTOUtrOjiHgbIZXx5OS3xdAeEU1xGBnCjruvAO+IWuQHbwbocOJ4iA
5Kb7ebz8d4yoktqRtDn+575iqSMSLS6SvG5Rf4TjYSRKcnjdNnLgYXQehCy/8ECmXcZuCBJJHOH5
KrHamy5lR1fUbpQ+Rz3guY1rZFYH0xz309jcR4CvqTj1OpASAMmBS944JL/nGj4GIsv4skK/wtjf
1Qp+vK9seFeCT7k8iJoX+ASSKm/LX/2FWnj414L7MMUSToEJ+7aiJfJ/YJgSOhL46mwJIWjyXXQn
qwxi1ptsDxHSfkYph6EpPCOiwILqMNrG5xkZMGB41YyqyHAlgmHlrvXbR1NpYbM/D4vfn52a4JRC
kkB6FYlRSFZAUbZh79pM0x3yg/9oj3UYpFzbdu8aSpGc97i4sD0LLZKfMuOiwjrbHbdrREcETuh8
b42q+H2WFjhalAa++Rtqx/Mah3NV7fr8OSDJSHYXnjDBcsKIkRss9pl/ZM3x09qPtAhaGMCzRfVr
+6+ATLkPREDnGrnSsRWcveNV1QJHbc4xsZ3HxFg2SodEn2pOuSCuf1USP1dIr5yomGL82Pmom4j1
H/hN3/qzhWURbdlpxIngGxrvk95Y90N3+crTSjCI0sSnl6gWcXJtsFhZfd0Sqqm3uP2AST/7/F7X
7uOXCIv9NZRu9IAhxTTn6ht1nCWFumLpL5SE+YxPUxOw6ie32tRa6TCW/wMQOHuMLJk8bIB4n41a
7TS9IhxE7QNWmFV037RMvX+M5kk25P/P2dHorYw8m0DbvD6ASSbTl5xteGcHMUINk6aKgb1CgMtb
y3fnBv6/HROAAG9YBb7lpk6XHFiKk9Avzz2udw4gAu3KSjCDPgKVAS1OH8BUOzA9GmeIeAcxGFIo
h1Ify6uXaXlEGhsUmpM3K0W7vOL0EX+FXbZ92gDuaX3pF8oFKWJell0qMsaB8cBEZcG643G+8StW
x+29GaQKB1RTJH3CHDbu7FK1TBI/uKLOzhweSDr+M5Zf2t1EO77JJr4U3kIkhqGxhtaGzUPl8OkO
N7PzZmyuiLmGhcuqUHAT4SsfYEUlwO9oKHR2qn+28HmMvFGriVE/phC3bG+Th/FIFe02Xtkovl+s
aq1hWMgNdY0blsK/Votnxx7xPcUWpS7jiBI90UnaII/lRL1PRZ4qp8O+g4+gnOqAyQTj1SnBEYm7
tkjCwr64P4vI4LKs6zNo3G4IV1bxEwXyPtKN7Evqj9oxobtAaxz3llRS343Ot2yyQYQkPQbII7Sh
OG1LzBjEzjV9j60D9T1TnKk/+5lTLprFCjRwEPKwVUYcX8miiwpDYpCMSTiJG4o1kFJ5UthcW/ne
T2Urkpq1ZlebAZ0Elqnpn6dlDBUP+a1jfUX8kyjcVgYCMIUIBQFoy2d7gDWsBUC71gXJ5U2Txwir
OyfzFFHoUxriElh5R8SejVtbgh6ELMAFVFlaBKYljdOIHUVRaE3FtRJMzZ1jC3JyQZ5zsCirFrxg
FyuDsit4iPlk8sJGP1NTkw8rCZLTSrjjeyOGkhW5ugpI+zCzuDyXmrQ8FxaSDteG9YnvYA2jcsaG
+usxlemI2zrlfcEyBm0BsvPiNyeEhW6oFN8RJ6yMJVX8FebhKJWQ75zPIsPLIo9f52HtGg52HF31
PpIyqsb8sJrbkKMtfq3buLKgGS05ulOMcSWyjemRbboiT02csAVabH9N0Ln+z+O+1N+lW//TXqpO
fl+5DC1U3Dn08A6oLKwF7TvQDkKlLVmZPu5f6asmi5anbQ4tuVEDFtYsUdZhidxpqIzjNO7fIcff
yQVCwT0wvP3mmS0YUOpIzdrbK4ejDqvPc7d0bLk6Sk6bMvLGS+U4i9scsA+uwwMH68uTQ0Ku6yV3
KQjdBJ/znqjAUIw82rtRQZXxtFOmY2Fq3pQHlVKyIq36s39FPTOUihu22bAe5GuZJoG7HF+Lem3U
EGavPG9j2rpOC3fdCL3/vmmAFxKj1eyqcEEGSfFyUK5XckZq4CDq17IqC7gjUPZ1kOaFJg7BHm88
arwn71CiF7Prxit3A4tRUS+PjTBBctkBTcJ2yR00ZokN9GfgRf6immZD7HnqU+SfO68/ewDxcxXA
Wn9AnzrFZECutyljzTLElX1N+57vGwlBCoIYzxigI2XOqChZKDtKq8YKEgPsb90GPEJ0uYLNZZb8
AsHkh5hFiDKnHEZ3JfM+WuVcz195Imeddqnl5d+u92wmRgPLVzuYxhoJvMu82UWumn7WPDnSqS1A
ddIFxuO07XLRSxWaj5CS3DnKSg6jREKihSAdl+sRWa1pIzp4AaGj25VdKVoeGmVALb8MR7JEn95I
oZgWfypX1hz/sPf3bVoorLFZZFztvlWf2Adsk3seTJv425J7mVYwEtpXQAAjmJfe9f3EPdweprPS
kGpXRfMiivemJusQZ4CoHk775RuPrkmJO6lnszRriYPV1O2lN5wf1xKtraM/sKrcjiZw0yrxErqe
YRt8Sav6MciIFqe9K+IvlnfjZSxw+HDZ5EBlybZR613E3nzADch0Y4NGsv1WTf3gkeJN8AxTtPci
AWYMcN6Dot8aK5hgAHNiJdlq86Bou2NyXHiNy8NAt2Frb1kNSNUss/TxSoOUVf9IYt54tSWVhz9S
qz+elwK/o5CBoS7cMC6Ta3VT/UjUKy34I7+7sMfrRMzOZPsBSaa2Z2Ax/4VEJn8K1YHMq8XD0Soo
oYzqgjk0m0c9R7iz+9K5s37QSDAJu+Lk2jO9oT8DriB0GfhQ9FPHUgBnsHda0WuI/3EcpaInVZhz
zVUyoEGbM9V/yt+j5cG7GDfJp1ruW2/C6DoyM3b9xKvYdB4cXuejsLgx63cIl8LcKkxi6MqERiYX
hzTFct3/EohpVjFA2sp1CJofxBqiZpYK9aqunyQOotBl+zmslEcK21j7B8289YHS0Xiw6dQAM9We
x4+I/rp6/0mQum35mGsOJm7668n+S9WFHYaQd4YcZUyjKif65punIZpJfVYbwdujb5XHHq0qAVyf
iKB2sNcKQH8vBr5VKgUlD6DWc6vSFw1s1MdRgYBOBDqoNpKrS4aHdBY92+5Q1jBn462Lzm8ss6UU
PNntvSyJwlDeoxQAn86NiZFlWd9b60UfkYYgdYxpGW0k+JJdT0Ghu8nXNc4eHdKZvMcLphb9yzVR
s1lx0ZEHIURMo5mignFRAU1d1cVnjyefw46tq3dte/3RsSjy3P/+hdaOMrGB9AmaKl4FF+JMxavm
HkXTA8Yt6cYKTR3FVhJSWUIrMkCaS18l01t5oE6WDCFtpy2dRlJTisw6JPJ9OYuiHzpWZg4PG9Nr
nWWXa+gdMDB6hObn8o4I5zcYDdfVfjJPf1toWqJA1wxkjblj6Zh7LTuRi8qtP6RGSOMm4f24qPAJ
GS+WTqSVoDVNrwRopRrktSOvy4NtFP0okK6wf97Gx1p+XhDi3SNihtO0UNioHu2Tt2nw6nDzRblI
7ziYWE8i4WwKvVM7QNb+R4MvMRZ0AVT65ZY+L54fUEOYr8/pD2r+JlUbNNgVZ3VJztwUd8YfCMU6
HZTxEh5xJyRy6cMCHAy4PShPiSrmXr2Tdldk12WVAAe5ktF4xwLb6S/lDT9rPmHm8x9uDEZ1J5nD
4y7t6MuTruBFD7UPYpjuexdoTtrQ6yGr7p45BJyLIIaq+J33oZ6N2bkrOkr5u9qKC7MfnWPIKpuT
SOiFtquCBAH/kjz+cSnL8avD7xEexqDmS5qkVB9C2Mxu9AzVMcro2BX2eTmvNlW7NUWG9+XArkoJ
dVYX5wt4HyigI//NWjN0/629/v9SQ1A5IXkMryvbl+zkwxif21wtdB2jb7iM2XeC4nIsC8ovWX/q
8BwNFBrS4Aq+R1MJpHBcsYew23wkpPZrQ47dWHic0brcYVf9msGyj7kdByxSDfy4f0dPvP8ueX3O
vNmZ9JITQEgIhMLRQxRUUnYTL+VSY9kiRyCCTAP25y3vqwPHUoXJ76qTwsvj2Fj3l0Nd2fa5kGG6
5YD5wOIEnIwh/RYV+AyHnBoOdlMq3BnuKxOYP2SA7nIuo17tveKiQGXEExrlTzdqaOLp6n3WB7J8
ssxRid0flw8xCg2EhW+HpSRv5AEGAsGzTpzgV/4wc5OPEQvS40Cv1D15XviQyJX9ZEDEzvKu1GBJ
rH3RKXHvOshQzeZ6cRAE9PJXIQxF6czaNO56FRDDgbMIhgOvP73HrEBEGVodn3lcumKvLoSDoAde
PVjnNyNJb4gAoESVYaJfiHTfYwV95q2FP/A3GDSd3lVitwWHwtRhm6glBt8Ow72Ylze/PB2Frk4t
YZ6w/lFuoMBbzD9yAQw7GKFmzT703hNaoEhC4cQsJKiqpDPXNXg09qSzu+Z6ljyYvpdVrLayDzpZ
kMPMgsnMsWqmaSQ2Jp8KXd7e1q8FqMxcu+veeA6+YaIFMEabvxMk5ln20n0SiZGFuoj8o1/P/yWU
FgsLu0vSNGAncPl4RXiHr+95SdWJHqCQUK191H65CgucuAdFcMl72jkdUhPG+cq+mJmdy7UZ7NBN
WM6tGobwsbeeLZfhlMWL7DrLiqeDP+K+ENH7KzRS0nueZ9it83awzMkMSI9K3AHl1qd4lNbbREUi
Nh3NaOX2Tlh+r4cOicwdI+N5jaL6SeZBElGoMH23JKXLc8zxQP1lKxa+ITwn1nmZF+0LTU78pdw7
kZcnO8ZIB6r8YTnqMzDvEID8H0iSjWy86C6I+LitrKLNe7ntySPT2BcruzC3cYNJS1wlOm5yX6ie
UX2aCLhOHbUypj1s4HQuSUqkazG7peGR/GO4BQoQsxYA/coJjQgphtQi11UYkh2PiSRJzu0yjhVg
Ca3snbvchUBAki/CrUM9XREHIHkrtRlaTh02pHsrRxpX10WgphimsOzXVl/e7A+KN3x60p/I1Xgr
nEj0IV5gla6ePijrHWyEpIZWJnlxT2Hy6pwHJJoc94YVWgKJVC2FJQtUBQrR03pHNX///FP5YXVo
CpIloQWc0/Pk77XdQVOCxnwapJzCf/0cG5gEs/Z0VR+Ngrr6zJgb5SUu+7eXgGcfev34QvwEY8vw
g2VTprIDWpryAAnmIOFC/bTZivbFNYwHbATEP1j1EYo+//bHZ4q9s/nQu94bGcsbEB0qIZ7vxD07
D9VtWwhsCbCLyr6El6d6VoDUu8m4l1nTeYG1WF10xtB69IywV4I0EG19Uj61ghfW1aiHeK6G6jm0
i8MmIL/42R0GlsvbOfJ7wSvnCkNOsT7Cvjax944jSFUBCf2RKWxvOK2eS8D55ccdPbCLGBq9xVNL
3LVxk0NfA6/IuNDyq+xhgVoC0NqdnS4LskTFknO+r8+4U5L7u8QY54gYoaZ49NXJgm2vY2KUZveJ
Qxlphi2b+PXLASeaJdHVLlQ36siu/hddRj2+rMOpf5tGz9h8wf6tXl5ILT2KUzTrBvIXQpVRYofX
k3YIX3XDxzeyNZc9T3HTYRejN0b3ocMttuX+/WFF61qPkzEcU4oY8W7uBK0PFz0GOhi6KlPq11MP
ZGtvmBAC8DBkz/Eaw6qzfqrZh+y822f239IrMPbJrLaCCvW6NmlFLHZlcRJkZaVfkHmHtWkBwhyu
EEc8qZUpJRtLBcwtgBMcV1Jibtv281c1TtJZNVtbmzkE4bexAecZZeEBUzttt6LQ2my2Pv5/X7y6
nwlgnxIJpm0wDha4Kg3RTz4RtyCM/4TY12m9TXvl8fTx5U2eikNY15Prw3Whc0j1BmJ/eckho3VO
BgRMAfD5FG7a1NnA21nLOj+Yn53UrfzKpGDE1f8lSMe+CwFn7XB+9JLM9ErFY0zFU/X0oJlvABaQ
4m8oa5EgqZ6RzyvBQ+pFcL9d7lUrOPtaXm+vc+1fc07qqGwaBKfo+2aQGY4PdfnDqhVHrqYZC1Rd
5diPmuENbgkW8YXH/wXrRqextnFnB+ZpYhQf7Hey5dM8isiw/4/PP68d6abBnVqRv9NRmO/8tFXa
TJmlNGNIyXmA9ncyOLzBcbi0zxcNIKVuaoPeZjZEzx7cJ1BML6YqfPfLDzT2Ak3V9eoRudjt4AUv
TNhMDhixJwdIAKYrgqlbCCf1op2HxLI2qxwK0tLmcF0dS0ZP4btS8qMS4BvLkLhMfZvUOLT1xXTn
6Ul/2JJjKTqiRYYLSDfoFenYmydxtd/8hSBIP2Dc/g6oTVj0zHTooueAofcVmq6lCrXS+rNH0TiH
Aq14Sbw3tnqejfArAmzy1u7zcwwd5MV4p//HkbFjJTCagDIQ2Iozh97c7xSfy1VjClY2wSDro1VW
sPhtiLD4H463uGGmP87DiweAwI4JQIOh4g9ZGIuMgw78q6smjw7yggnjFN7QKJriqOFiennWduy5
Fe4ih06XNQWipst6Kr9QV2Yqr3AV1GMuw+mkvN7h7sb2DZtMaNvWrkRoFx85N0Q4ltz68DmbXi1h
mltWJ3WFu/cdfsfACQXddpk/CGg3fNLoP/ZeFmUNGjp85MjEXfW8IODLbyAi1EhZRZ82Db/3Sg0M
BtGOGQGIViGsPv5kBvZmxjk/KeuTzURLZ0AtqhqrXtfOEHWG/+FS8IpFlJs5R4x8/bWm+wf4qnLa
LcK5+tS7VXKasHhNnhyPnJERVYMG5g/vcC+/y+bQKAkq9Yhu9nTAZQn0QS2RVguJzCGBphKXtfCm
VfkutmCWP21iX9oM5mABzuC6YC/J4DMbllAAI7r5F2JW9W8VU6dBp4glqylGGzS2ZWRCHt41EjkD
aO7WDXIztuMwz4HA2ulvk2KCvj5kuiCLwIDFj96ufYsm0ABQ+qnkClPEsUYpUsz5H/d+4Ttb3SeN
IbZ74i/kbpoUF0T7S6a/GKngMn5k8ijwg9yIHH7xo2fuCvLQ/AXPKuysGF/rQdWhLAHX7wfboQTX
/FCf7UvD/hqszm2Xny2EaDlLaNlI7zPVB4u0GRFvraLKu+Qwt21T6jrqKkwjHq+280KfsNMVjlvl
eAHLbmnuGX/R6IRmMRdG1op/tUVZAuoL2xLzVslHfIB5qaLIFiw3kVEifNiWqthWd0WcQNuWaScl
SL/jX+/vaKwhJNvPlSGmWcmgpBPOJ8Py209K7xXH2eIpD4DnDJ4FWnTnGwkxFyUf0Knv9HHiatUY
9eJA2IcaOXccwYwRmJUk9HZRIan1vOQ0pI8gMTcfKTQMVjxngdfrQDTsmNavVBFpjMGQBwHl9CaK
2wh+l+mkDI4TINtKBlMtb03gH/XDRaMsRsPq/snIny/yL4c7LQAlSq0xi4qQZRMpOlxcmo6lxSmo
z/tqyXHbh3wtZm6SZlLycgpdG7SO9s+i3VehQxR0+mfL/PvZCoN3wQRXJcEdlf/YBmNQD0IjwIz0
VeiVx3OZjNfsC7lpgr2thUXAUFoPJBp81kntQP09a/BZ9Dr12ZCJ7fvB89FtMsRLC2MCrFcLty6w
QdbWIjGR9+3PCnxtea/ye3CzFDc3cS+Lbho65c9IOrIJEUvCkovTonh8oHit+BHgHmt6DuP49tJP
wHQymlXqsyV+XWsYC4LEUu3Waxn+AwzVRtl9kbHNKxAf3dmaqZIiwOO1Ox3QQrDCKLqZJOiPgS75
pc4DpLrA5JelksaJLXIDbkMQBL1TqQu5n9sKcZyvFLeMLdxLSGC6Etah5FLjP4Qy9ZYwl3kr9U0a
VHWKNxr0Z0mR33pRxTrR+id0okIbjXLp5VQoDpyFA3BRcc3eahW/2sox1O/Fa4RjdrXlW96sPVuG
iHMgds5SrqgQ4wPSB3fQrdbzi93CZnCFqwat9p9orD9e00C+b21F2C9/vxsc/mVstUXnPYIKovhU
U43h3RGsBvNrDF8yAPOajKLwSGvyFCS+CVHNxudcFsxvH2wexIxDXMfwBZLMosnW39siIIOOODyH
c1mz19VBP3vwoXtRmWyzJgozE6spX8Z7z1EpK5svT0bTLCWkNZY6NQfupsmJEUUfEoyZF0z9jRhG
a+TajaM4xuR3v6cZv3lRmZvGDIZlrEA1YsdxuoxsYZaMVr6Eux7OlKMpu+CmKAPzdKpAyO3ExOfb
kyoZc8LtaqwS0ogumqlgU36VrPFUC7UB2ozHvYaBUYWiHers03pSk7H7ojfP4j/blfs6kqndDnsP
Q0Qn0bQRnCGCsONUT96V4piBl1S3UVqARhIyeD9B+NBUiYtnrUyNJjb2Bg5uQfsJKbU91+gb7Aw+
zgZoSzDh1GPfVSrrZ7toglwm4KPVCo2FupJcXl+ZXW1Ob+P8qm2vaICZ/kVwT3Vlat+8DfTUpL5X
gEEhlpisxD4VISArU98ltuNSLTMkOKquxb4tWU77Sa6GfxkqrcgRSPZTAKCHuPrL7VRVFbu0qnzp
8/ArlDKLC01XxEF1+ApGJl0ngoH3d1V9EFi7R2CHu33cNdwhUKr289TbpiZxNXgTkwHKztafB8se
uYNH/wGdDYEImhwGGUlYgN+nQRKoKTvT9MYP8s3lFC4YdGJ78s1su5pkoQBzloh6RjrXqjIhqGuf
gNck0xJnaOg1jSI5XnOc8Ucg1erw7Y3GKvEB7unGmgQ50LV49vIpKFwHcxzmXIfMb2YbGKSz/CgN
B9LojdKL3M8F3kJtCYa7DUj6mqfE6VZdjS/Y2C+YGZwOkS+QSBHc6Nr+LK0roclIXNy7GCJ9jPzd
umkDY3yJ8WCbGyu62y+mibsJi6giyV7oyy8ZpySnNNEp6V36UF6Q1cSwrEeBpXFkZSOPZp+diADO
ocnJVbjy6P4m1x7gpAms/T7BXWbEUGuj21DTTnuYS90vsAiqYF7gIw5QBL1ipWVeIhtgzoLeuhP2
/irODbbVR3kuFO6a1xuFlUg2Uxr5st+LuGLsgbzXL5vGzv7FT7EoW8D9I9X3dbZwyuWFUzS0QDTF
RiEk84jwjiiZ//i2cwzyD5N3e45CbVH/GQKHKULTeIVEsF8Suaz7IgZ0pF2a0ktjl6OZpHAVkOUS
UDXN/W+0hD4l/w7+ID6jMMG7UzKpQzH4S9azDd/GL2hIcCfrZ/ven5xiTFr2BUrdDFO0MizC7Q2b
eD1wUvLRNm220x+5N4rd5qMI1KVu2e44UfgHpiwJefGh4RthLygCWuztoyPSfdtI2PSKkE1gyHwS
p4mkYmjt/LJwiRaQHLtL2isGo51+lm6RZ43C878dnd1H7c1m6BnDD9lw+erEINHgs+TtjynGa+c7
k8349i86PbyaipZDWlmRdEfI3nEHFa/quN7G+lcRiAhgM3fEfTaVG0N/d1NlfbXVN4ISY/dVH3zQ
0tEfTvtpXBcKF5jX3ewST7eyDm2YN9mo9dHl2yEfHrQCsspJUocC2y0MpXJlOldQ+gDA2GZ0hOSq
2YxTEo0bJ5nuHpyAv7AzzVbRl3WdXePXsTvg9zjbBMMtEvZJq+ZFlKSb4NlDDN/jpL6g9yWpexpS
hCYaGTsSqW+/UcBKTBw1qnHZdulV8qDsamC7swDgr/YcRAfZMiiYwYAwLMe1pYodMY6cFymeCJwu
Xjwc3D9MTGsZpHjP0PyuiS6Md5rKRit9nL5/oM8dWp1gYRUFQzlcm09j3axnBw2USeHjiqM8Tif/
VpDStOymsdEHOKrxRCfKjjRumns+HUE54NegVpl/orb9iQvOVaTDL1KrCLwMPK12jvUGAgYVW/Tj
Z7DCw3oJXPE0z+GgB73dap2COvjWvFWXOk7BfcGQri//VeJvolUZ/dFTGnDfq4ziDAY2AsjU+uXY
YnCmH0e0WT7l766ZyRfIAAk7iwngi3Rwxb+UvtIYKJ4+KZB6//+rrkxIc0Jdy5dEc7XiQ/N1D+N5
m7Yve1L61A2Wz5B67uthUtX6xTBpMdaUb87uGNEgIAUXxp/6Vfdl+MHDIyTuSObg0cC2SpZko3Em
gPDT2HvoXBKbHh+mxuiYLPhpirHoT9H0TaiPiRYqkN9cCousiG7zpjmjzcuSJOn2wXQ9z85xG3xr
wZ4RX3VYSpVELxK4PN9zjGmI3Mp4woQUuzSqgKXbJtCogis0ZtuhcHmolphm+b2MgyGAgN0a+xwJ
JF9ysrM6Wj5X4wy7ED1QvUqzb4PdHeAlQqiqKJQW6jA2H17mjSibpJjmJE7eYeQTeZFrUbF7Di+y
URjxpIxL3vokxCjUJ8z3UUCL78nNcXtWFIXdI5FnVAojHjm9sUsroTqBZtB4kqu3Gfhy2Mhpv30s
yCLQ1WkAyM6uVyQmpRYYjZv7elVFl89vCPfl+zIHZYh435lyo9MHwxuWqOVDKO2EJlglPx9+Kcqs
CkD7TNYYERcLv2xGuuEcYMy4vPmAznF+TuC3lifC2znd8F+H0BKwMr9M9enriH/kw7ZnmxmOCSl8
1cGoHigKNtfqKkKKtk5Pkn2XnI6JivCjo8oBTvg2pjL3xUXs0rjABDhV/cH7gY+Q9fUqKz9DZAGt
Q6OI3WBFbKft++9FRxxsX4/QF3IsJ30K9GudWS7/UL/EH72wmcOcVNaqd9tDBalBoVjFthPFB386
E781CPTW6d/W0hXG4x1jDuUnOm3t5AZfC5VcZuLpXPIOeayl0XHyZhidDV+Pygme3ttCpS0OQl0B
P0wAcwbzuiUX0Axdrghlx+2HkiNwzk3xu6J1gQeL6ByChUJISz6FTT6Rb1ZnL9fgAq1BLYa2J8ai
ky9pcBbdmp/cGnEwdv+elNPP3OgHRthn14oMhdXn6NoXQKVaum7T2xtKCgi5q1vds3Tv9LnyM1rT
MufRxcQXtx1bJnZ78A6ohoZlx/QNWvv1mxV1bzoMt6/M85yHvh1LMmCGxG75yA2a0wo1IbGK6o8L
F5u8OMsh8oMgfOnZaaNeLkE9vASyMmCz88xKtZfDe66HWvYVn2JkwD8kj6QzKM0RIep4+KC3b1Wc
Lpn/Li6P694yn5TZvzUGTdeNK9rm07tsOs3i91Zs+TCJqzfH3SG1b0K2hcFnQ1F2sJCGxO7NTOV8
jZoGlCzPUu8RQM6ruKF0ZVrWsfbaN/ksHovQUnz6aOXGqzSob9AFaFMRkbkREdLXBaUsmOSOi6Qi
d9TIM9ggt2onZml3IlbUAANRD9sxBeylMzCqdV+E9b/z0gydF8uMuVNgZRQFTZ6ovI10Op/G/wVV
LGR0J4t58bxzz1DlvmX6L7bY2ykH692Iak2QS6I6C5sqW66PYNv/YbrQSBySck5zvLYwmmlzYFC5
J7gWKCMMPUeUS/V4rkLvXwe47rBlypv3dGJIvyfhPrrbRCP72e3wzIluUStr0UJMwOJB/bvyG/M6
ETM+RSTnUgwAvqSbDlfXg8lxv+DXVl8JOB2BTHT2v2oBJfE1miy8GTGz9aEaLmLC9N/NB4a81jJb
ymcru+HfyMH0C91rSmV8SBu2XY367KcOC2pk5dcNR9P+3TxgHlgEinToEa4QGOZ3gu/5/PYC9J3Q
dxCdiVxxAh86fSndhDANGk5M+PNaTV1h/izVNlr9eErumWZyMTHv4YJjYohm0Lnr8BqmdP1WxxwI
ywr1NvSryUOcALvpeG26t9XzIBeG2tEkiax62HP1Nds3rzINidv7ZovGvM76xSFdZ+7qv5plVyBN
iep4M+R2bj6Cn2E8OiBkcqwIBLjQ8q7Vfcn6JFblrMairMlF9en51ZaR4RY13DZN7d2R9Vwo18cY
dgyul6KpdirL4+y5xijLY6kZsuc0u1qdCaTfw/xV+SvH1uGzvE/0Bypg1DRnP58LQB2NMZMA1X0t
lLF8DcwWpUlNWas3alhAz95atqA17KlzgasikiVWbw+qrUM1/k1BVmVvTvcyQ+SaExyNP8bdUYx1
D6sOgVobwriWNtjA/elhqlnx+Eh8Jjpjg+XjlH1IvdXASYp3zz4Qz4qMBzoC0t6cQS/ehXHitrYI
LK1Az+LKUij+UGUeohjQY6o3JHL2x7b5oza7Fn56W/qBU3e4EgSl6ZX22hgrEvQx7m3h5nNGqn5g
4KIG0WjrcuOg2B75Ul8JEH3Yxu8U1orac+IV8/DEbEp7diTVbS1UYgE8c23em02DoHV/TPCBJexD
CeJxh+Yyko94w07TCMjpT+fja8L01yoYLpjeDQj76uMmGBpOiny+EcsFJi0enMyoNmk5VklvHFRZ
X4feFQO+8vHpf/AGo0Oq6bSg6dIAyDiDZ39g2uXI5g+bMNHFLnc94ycbzqpOEUJy1X3O0/TujBRm
aHddClMNdPcslaMdP42rq7p1umu0fdVzvDyB6J0j7xLlUv8lDQseceTxtf4lc3LgDUi80TbK/Mvl
cNEcDri66QW/oPVfaP9XmpM8v9ImauMS6UinvmS5M9Kg8Jrbkx2AbD6QD0aQhzyUqmk2eVThPpLr
Np649NWAXr0gurzMMcU+C39xyc2+mbJtdr1EPFidyxPTE5iuboGut+wSmJIQBylFUiHt6+0muN8l
F+WFgHLmL1LMnRNqZPUU9oW96JnBOaJ/QX4HHoNNxxoeyWzOOmPVMqPvFfnWCqfUj1cJyZ3RUbG5
lC5XiVa1zkDxYVF9agPUMBYiMPmd2ZoZFl/h19m1283sYvnlZZ0xJe9ckw+9A9Wu4myULcWEmjPp
IfkJdz/nzMviuPr4nAAEHCI20ae0a93Qu8cHY1NhIH6k39hPgDjJelPu+LGcqFnhmc2UW5fboJmp
ZeXFOJOLIHBswbwKWwmmZIwb7DY+MnTUsicWQmSwVPZXFFEqfkgltc7ssd9NNEUfTkmCN9aeP88T
ol7NwS8q3yDtu+pbk1AAT5OEm6FMT/m6r07wK1mCK9sLSbCtqf2doWjgs5SGIZ+H1VfW7vVzA0Y2
4HYqk9d8z84KWC9yYnBsBUNHyIljZTuO8GrYzPZRrX58d/mqMfP9EdX0DHGV23nxqQakIW822fjH
2y8FegQI1+cn05aoCmGpPVWySFS64YNzQBzTzKpiiQ0QeBcr9wFMxeadH/rQ+zG/XwS4tUUneUnF
/qP+doGgbl7afrmJjrWORcgHc3TaN0WhN2ZUi0ldlRwIfyCNN9v+VSO0E3CVLJyhqMIK83CoFLXW
I/fTfRXOMAy5O1jCq8RmKimw0SYThlFp/cbK6YWPtevJCatq84SxEvugQPh60/jSMgURHXZUjOrl
jF1b5qIfi+tyk2f4/LUzp2K2dT0SEGPJ6noGpdi6KTBN4yDa/WSWF2RwIyEkCGbO6oLkN9nl+T50
WwNFCQpSm2SvFXovvC+/yd7DhMU0XGxL+0fm1tqxIwFVcQyQ1lrtygZ+9Az2iRKrIe6BNUvr2PB4
TltX7KV3s/H6ENASb/AOVv30oQ0ia01RNoiigjpuJneKcSGHeRr6hgcAwJBoh01QFBRgv6Tmfytg
IzG2iDmq4qIhmg7krLY1uV+tmER0Hkf7JI3OEgJKGQk/7ar/K8D043AGjt7tB8lRQ/Ywm2QHjZD+
6K3Iir18zfmxJbeji3b2UhrSeL0axkFbRVxykKaggWTJiiKvkR1hbhz/Rj2SMfrIeFN/qAlPoaLW
BiNYqUbEXaZAOAJ/QHHXJUlOymHcnNjPipzktl+YTh6sKSzWqBS+qStR1CuYxfc7C1LP2LI5KSPw
4U0rxS2lk4P9I61G47odwSQNVDpZF6xNQHsYh8PatrEApzjU7oUz1nkggstnJs7MrAXYlQaxQy9P
8sHNv369a2FFDBadsyqAC8qy1iy4iu+EFHOdULMGLmm56Vj6biX3SqYXzkkeS1f1AnMn0dHMw9/b
XIYOo9hXma90rQourdfs9XogJMdhijbgQXeHQq/QDG2D8HGjo6QW6NhlacrHY0Ovdv+e5tIeQnxp
lrVWK1JQcoNmMsHaPMat0Ugy8iwD5UPeRtuTMQb27FNfzxCi8pIwk4gdBgKPxfPGcl4JSV0BEAhD
GoTGuZErur6FCmA4ploPwcixo8Kc8rSVbalk6qm1Z/7jOw4dU4iDkIcbS50vd4SYSLK6zDZ3JSMR
lypVEeQQm3tGortwcJzm4Eo7JrOGRlp9+68d1uNfk7EV8w098b9l+5oO5hnzaXh7uL5PjOkXxKxK
qIM+tZTSSlc6P9b1U1SXmixGpZlwKqn2gN7ufsuUAwjE4o0grNX+RuCCrooxxx256DT3sloOX5vD
X8Gz36dkCm1N0f/fWh89F78SmtJDSObsQ40IGJDx9x+4uFGa2VoOtDmOtNTIgKzo5hQtvSwXI6K3
uIGQWVBXpBb0q3VArfj8MWr1JtlJShqVALO/lUMljTXkh4n4BlyUjGRJwR2ox1ZfKELQwwY5lXLw
AY5LqWC/+M1zVNnsWg+AI61NgUpYxHQ5ir/YBvc7lcOIljD0YNM8RQWFSyqdK45b07g25aUF7adC
NVBA/xbpO3XHHmuqxQBJlwK/rS7If5CvFIEAxQRRsSXGoyZ11h0yeCHE7NmdkXxxUtp+AJZqxchr
247JHVKjmXk79Kyad5ECDMZHSHDmjLiXoyXPAN3p/LvWTjU27/xDoERVJA7ybz27rtKZzm9xAXP8
/GCpZJfNqJYVw+lPgMqG0dMoeXJZpQ6WrPYqNuc5PcgGptGav3mqqhRSlKXNtFwDbDxfGI/7HuF5
cRyNth42L4jHyIjj0An6TqbVlpwmJ5U2XmFKoP4jnZqFT3NXDKF35x58veLMqUXL8Pm0s/vpyNTl
BlJXYbNtqa8eR4FKJZMCwXWYoI7S8zYdj85pP19tVAMSJVjzgb2XFWTKT/mkh3GdPFLGyxNS+i5x
5xx7gMxokb8+Q1eKfqef37uwgopyD0/MCj5YYGAxS6ECeI3clU2KRCHSsu7TarjOjuYhsiav+hfU
1TekVPyaH24l/hHX6jPoRlSiIHfdgE09GX+RMFacVLTSQXcGJMdlEA71BBq9I3Pk5U4YY0cBBbxA
AO7zDITWsf/R8T6eMIaDLRflsGVyFqRjCfIM5GtD7QrrcLk4U7eqjJBUcVkFpS6kYKdZNY0u4HzX
fWOQLSj/D/9dOVaFIA5jv201iMZ23rUGdjku4AnH9P/CGFe6qkj6orMgq4VVxwFJXYFEmKbUKMEN
QUzO/oq9jJ9dfbh5ap3+INTJXqVUZc+jZK5sJSAwz60ZrK8GaUwVZD0+g1ttdhqAtGTVIfLEKjpy
qIKj3snqBUstFI1uPSCCkJCnSo4kDVbpprN7FN1X0JRmGD9jzJWpCIGcbTrb6uZwiEvWf67gasI9
BgFDcRr/hBQ6Uwvrb9NWzj/zs/ggFfyeD+QLjAynen8erPpnCP3uWzEE11Typ8YG88D02m0FTTUG
YSLMEZTtnCwMSvWy90I7OAr3xVDyjPL4CFha5/WBgTOTogB4cm/2n1XtIERle+wSOOynM/sgcd20
VuNljRiRM4iyah3/H1caL54fEoiBmfglIbKcFa2YmmKgC2uxBLXzFjUXFjVg+YYMqkFdqKl4n3Ld
fs+zhki//s9hR8CnfK1iiqaLxisARus6v+G7h3ZbfFjPK3I+mXxTQGsUWuon6vNeWhDbr4yc1mKd
/eM/8MV59C/CwMaZGgJroLaxYJeL/DdBOokAhfeote68+gSwS9cyKhyxCNQQac6gElnNmyZgKJdZ
D4BM2F+9/xxvMcyDQii8xxZJ/ma/T+mYYHH6m4uUy3pCKETvGoLbdcSxpzKCnWAoptnHT//Iabz4
IgMBGmzYrk6r2GUMaoxJW7OCtvy4TBdiF4CEMVMXK8qn+8hgfFxV2EfSCEYk0UUaWhJFQzpfp0UU
q+f10ypxmluw3MMQQWEIinTg7MEOpn5eo4o7XXE5NdsrqW/4PllzVlTatPtyLaE+zvWYzL3M4YL1
tKdKAc1KvlRfFH+81pRK8ebanx8m7wpwNAE82MtDYjZVZaKs0rVeP0wmeRgiRUvoCkO9lTGYY2C8
wPe2aQmb/hX0+WrISJeERUqqD4CDJViLuqw7kNcBw1IjlmEuzJdplbUI1pUSuMuiPXPKRvrttAhC
ohJpHhCED2cli79w5WDQireHYmI361l59nO+97uF8UjMYO8h0GFR+JK3MpkAkB5yOwGnelIf+v4g
rPIl2jubdfCPzD3rj5Kb3g8IyzvsWsDMsZShZdqpzBTT5/EC65KZzbcBFS87QgJyrMsYBwTS111r
ACH7TI4iMVDjZruJAUO4uPriNRSDiXjKSuM8A6FQH87QV7Z4tW8IjevDi5BRJhBPWlRjsxU5S2bx
3gkTyyhm+Du4OwXBW+FbEtKg750D0hheBR8xPlPvwlm76KtRCS4EpN/GLzCz7tBDLoO5kN093JJl
xan3BBoTFJg8InQscwsT4ccLwU20133+mJGGFnJhXi5YcihrtfwjQ/s1ZH/45g1FVXJ2RRRsqwIF
flxS/mboxNCm8jxUlk0CmIUU6XJBc8AMFZBGhFdekmcR+q+CnaUHno/a5KuzoqqDfE3zdteaDeyr
xRCy7ab+Rte72ZbnRxeax1SbHCA7PC4HgfVo9YyHreVqnYlf74LGKEpS8AHPBdMqPFKSQ/r0sp8N
s1OxuoZJlTAxE8WxSPq85FfqPDmG6vg+bquUvyQDjY9cOdzv7zubRZrtsE1e1Jxjkdzjs6esPzvh
nd/wvsINx0iLTLOyA07BuDqnPEFD9N9vJpC7qRfOaFiPr4C7y42MLNtY4SutiR7j2dpiEiT4Y4bR
CL+pi97wCsmnDLxgSF5esqO5vsTYsTX5+pAuXYz9A3yG1kfPzhiMJO/3nLHYLsciYPbsqhDFqB/Z
qJ32i/h5TCLz+xSzcCe5B9HO6xajTC2YMrrB5uVzrOipuIlbXX54k7iKjP98ZzZQiFHmg0pKpf3b
A/zalhjjzk6rZkWDfS3V8xqkRDSr3GPeTYbL6c0XRKSZdBwWCSoux28kDGLNe2oIwCgSf+9TpFcO
VSNilKDzDVOR0W8tc6KtwOUNMtFhICnbqnQSljENRocI9N9D4UWXgotEyKd5zQ6CofyBnc6vs2/1
dBid82P6GYq+QzHIz8pCG/uPDibdVbIdvuIE7VitOnl6MyrJMfG5itB25BkYpZ9LfnBn0FzFGslX
3viMO7afPsXFoRNifBC/3dFL1+RUrzQyacKAfZ0sAh9K04vmdxps1K+8vuf2n8PoWk0YcWGAzFs8
AO9gtn0CI2HqIUJjgtd9guW79wobZU2yuJQvcCsEYKS4aDINyvK105U/IKhO9ncrEJtwmx8SA4Vr
R8IFYB6fQ+GFn3msGEaaqXIlyHlHjy2fMJMLnNY3k1S4Ku1Y0AapYGneG6JMnChvOonSDkx8avEQ
CdPMeT5kjI1hZPsw6qYOwHILi7EiHIZkJapTzAmv/h3/eLrsDKb7h9vFBAYRvFxnDEGqvLR5PijY
KcnBLn9chI43gAJU7Wn/ZR3uY3PqyTx0S8MAWoRkALPMtj20Qu8UfoISDLRV1ZqFItwkXP6nrrcJ
R8crbBRCbdqvjZYtqN0610nV23i5I43je2qC2aUPMKh7V7SeyHVNuE3c0y2O8yZWWFBKm8+RhXEz
TmzlT6g8G6HhM/AZrIheyaYzy2QJ6sN4BaV/Buz5RZhZA2A55a5lqMWvqAJorXBlQHlMjjzTmHd2
Vjds3lhfqVBWxoxprDUQ5IhG58IYVKUvT9fsm1tSUDItqmEkHtEk7+6p8rv7f9Yl7cXLKOj49sGl
EDfmLwghKHAZ5y0I0yTxw9rFaOBr+kQ/jh4Rtyl24b4I2y2xQ5VHOJ4CUKU8tPxT9kMrH6xAW1zX
pLklQ8sLiWV/9yjCwLHtC7CsIq1WLVhCOjGqCXxcMq7yn0i3FpZaHh2wPOLX4Z6QOOSffYlmcWo+
SPXbP8iFE2EyKR5yBuI7HzmnuL8EPqAJNaT+2yLrL1ioDO4b2Pf3g/0jWXoEX8US13qQSuBRypRv
oaPT3ehmb6Z4nP/nUO0almuROzaPY7tK8EEpuiU4Q3N0EWoxNndU8YoSVZ9wsuaBZbOWTf9fx3Tm
U2yih43uFI4cbK8qedLbzM182cQZhf2+rxIpvULKr4Ip3aytJyscJvepbpNDPEJvF9ajgBGEzV2e
FjY+oBB+nEXz5ooibZBMxF5o7xPbIWFxzEtq68AZFXgtkWPeTgEuXLO5eE3CqdAuOhM2zhPAz79a
VDtaJ3zSk7Jtnni0TNMJ3nnaYP610dsnC4Y8yCvKJ1ZHWwIDj/KAB08JHBUBA48h8WcogWWJTvHE
TBR/7iSuHcrZrAHPbM87+z2tbOE6YOoKQt6K9nvqWpOG0eiC9PwkVzMNRHanKj0xUve5BOHh/r+K
KqvC77HO3OGAAqvaM645yl+yS8cpoU7NXNSPNin6+Rm6ypVLvxEsdMi566WXL/jMcoAOBV6Dd8zY
9ITloqOFLA8jZYrK6dm/HiWsGIXZuIsKI5d/DOcMkffQ0NF9S5dUkn9RHhFj0w/bXYCiigm1ejr/
bY5Kplwu+uR1C+nkmAkRSBWIs/9OFD9azhP1ZL1ZiwrwrAFbBolsldMafr9Ph7IIhBlX2rR6rbv0
zMuOYQx/QZ37Ry5OxpoJJJsRrETnCYSee2U0eecGrrnUESmgw9/dvqQtYMaDt9XKhYUkgzoNsS/G
0cntJNBSRXcs+ZNaL3dmFBuL/rg3XEcrx7fe0v3Gw8MEUakCz1lf87V4IilEb4ll+GRCYkdtDOYH
U4RrG5kAorTCR1Zjd7hFRujPpraU44HNqoE2yWFnRU982hRQFc9gof6UaIX89T3X/I+GjNnR/w1K
KjjccKjEE7wtwLyzJSU6kj0+2Po6AyWQypZLKazmV4CfsUS1pAYD0FsycbXadFWK1ai/+0iUDojB
weJgDB7P+EOr72Y4ry0AmzZbTfA8Qj7fcxEJwxi5F24OTTv/pBM4krMrFWsroGGy0NonKhIE986W
GdP6hJzkziAlMjupVXoJfilbE9PVghirk/dbXncrKLb1X5VbJ2zyuxThCqF6MkBb5iyx7r8axEz3
3cmnr8Cu3IdwHXSw5mRJwUhbvy8apq5kg7k7MPLtF3OtlMrE1n3OLE0eMyzqazWfJJKW2qrcwhTi
MQ01WbXFBvMewOxjlVTiuBY6YY9CgwkHjFFcmya/B8FfCiX7Gk4Olm4zTLb08O1XP0d1goZ/Kqfh
yYmhisbuBQMUMNF0LLDAE3mne3xLOmwuNXu6UXTWK2CZNz3O1hI4pQtvot0ytZbz0FwTP3J/vUwc
PIe204r3Qi7diXtnJVb+KsSFrdE8XwK7bf7Ux1LkGih3rp0FDzU3tveZ/gogZG5QFkCvEmBrKiq1
yrTj+QwSUXxVlnTlCMjEI0YdiegKU1rnlBDC2Pd+NMX3xmUda/077Qb92vaAwUtrg5elg4bZcxyx
U1AQS5x+zPcqku+7wasA4fHBv6LUQ2a78ME0nU/yP3r5a5t6e/ibE9SCXfg4dCM5SJBCtSUNfkoT
EHbcO7PlvgI+sDzZikk6UGCddIRmoBOF8XqR+vqhMwPTohlrH79Q6g3LJzdG23LLhADBFEPN+Rnr
8eULDpW1eyr1XmNQJOnp6JRTb6YJSIt7yxH9ZDlE2KI6KHiyftBvx6QcAJuvza+O/IE5JSEx5Sne
La06rF7u4cWk2fO50hZ9c/FiAg98Or5EaxS3Y2hG9V3ivzmg/lUJoo/I70l02CyZ1axc2jFhdcd6
9p7Y8CHmIAtVagah3FZ2e4Tl2ElNq70m1/fx4Kg4198GuV7a1kvQm9cdi8RN8hxTexTzAvc6Nq8P
J9RS6/aGaQlLKsnwGkC//m/cnCYgrgkK8NLOeasslwTm76AzeKvzKotRKGvuYwpJseR8sogZYLyH
3SbBojHuApU9f302Z+m0UZc37N0kIQC+wiM2HKBwPTAKfsCtIBT4ke+N1+Ygcxk5fMXAN0F91JcX
0byHvQWgWG95/clWPlmpowHl5Z3ICdJKqudP6yZ0y6V1PxCiwOVEDuKMnaJxZqub/EViVMIsGOW3
sdz7Mgb0PuVFhWSBF+FbNO2aP3XcrJFMXOZnQHVgQNKbsE2CBucYcY/tk0nlqW0iCgn5B4nbzLza
aRZ/52gN5OfrmNyHhgpku4a/GdgJMrr8DN5e5J/BlGfTdG6axVYk4/hTreoJwvyprWhtWgf+w/8j
lXa/IfeGJpD1bDCoxc0Ny96FG+1FJEAI7SGG5LQPJiB3q6aDSnFJ/vp0pCBcsfnopGNS7qqCxM+t
jvH7JngQBhouknX2CoAkZXFKOCksJ2ewgss0kG5e9eMfm5gRks1i7VVLJrRFCiO4TXCPa3YZ6Hzq
suzfOE2WSZtKtYX2appI5VtpKsVvsqmASMODp/sINWc3WU2vioZUDUFXtyOedSrM46Rvn1CwWgVk
fZSzFK0EYS3W3yhvsh+7WbmDxw438KQnh7yU4PrabxenRQl5Az6dfQoEIPGeec1cGKJ2TrQIhTex
+d58I8947GitBp3qd7zGoKGEUt1N3kTU4hRf7tZWYSGwK3Ng+1dg2dySTR0V6JDhb4gdxYX1ufQX
BLkqtTrw8mN3ViNamTzVHmXNwk/l6KdhkwN+mr57THmfQKq1BzkI0NBJygBuz2h/H7OvInj8gTOU
KH8d8iP+v80572OtYZJh0ZzZicyA/ZJUGaOQw6rlLXb+KMowxkNVOB5Mmb87xBpJY7t2Fvq2x5+9
UaqQ9y0VSstHiHxgH61o9xlv9CRqMU/9B0Hajlwf3rfjrQ3hqhQ2MLC6u/xwXRmIEmmhavm4VV/W
RYyMcFqhm7Mpgl4o3qE1I/IA9fjyy/cEAuLz/XA6RjSdtzX9axoLK/5WLkSBEP7Ty3wkqCnYGqt8
WD+/qFbSEMWmUZTXELxc857/OCaXQDtr4irLVt3vXkzCxtdTVvy3CD7uBqkgJqQ6sJl+eiiOnCEW
8b+JnmOtQ1FqZk7fSEe5WBAtC1jkMRXiHmf7Fir6f7NUw/ia9bQyJTW8EIqO9wSbmBIhACEqeNaJ
g630kTrbfr4NBRPe0cVpn8v4LADVtvthHsGWn7ghmPHhXCDwEHRNeGdqXS3lNfRqYZiw5hfUCN2z
4FUBGnI1VhfuWLCZOCUZhNqEaUL5TJIO0yp73wtVka4FFoTl3PMY2MdSJV+1fQU2uf3luzaL4LRX
QNrwp/dLpR4+I93WkJioDAz5Hta4A5oiV+h/SHuosDPZhuPvtrDAxuCkANgROJ7VitIws1xRzImH
y15BMlJgzom2hyPJciFit99DGV4phK4CHbmQ8EAe6QjAY4L4O8z6wjKxIRrY7PQEUMp4poyOi+rR
6c2waWTYC8XGoA4bA+hw/wVayVBupQD3V/NIkevCU+mqINheJPvTRU64lkSzoEv0Ju2ob8rXRe67
EMqFcS8CXazEFbZwg7ss+u4V0Movhy6gHOYxgHzQrI+X7D2XiKih1X77FjKdOWzI5GMVd7i6wHV0
qAWmOB5t3OuW6N6WjeAkoEufJDr/+Gb7tuQnEbmRmOo/sGG/fgZRczPsnFCYBZ0cV+iFacPDYZg7
HxrQ0Zfs7qPzkGwW97mLzRSgJugIosdOUVYXFBwoqjnuTfL0qML5USlsZj/8hZx8tXaQM4agaIj9
wAkHVnEUoplsbBrKgtG5DyN5LLTpsKK8P6SF1iz8fJvKECGLR2vh5cspAKjHB3Xs0kcLv7kM4pzE
6B8zFalBJe00Mq32PjT4aciEO8jbg3O4akZK2w/R2NJuyWF1l3p0MjK41mIp/qKbWCESI91L5HGc
sHHlcmdzCDAPAdJmiW+V4AjTn1PHfwgUgNq+zHolSoPv4RDGMGl6E4w65HonDwlDJJmdVW6yYG0n
gYSqgKuzoYKnPmIqXSDhnI2rb6cNV9H6GUaeSoIjSOKVwlBSBeqr9aq/A5PESwwJqt2x6M/Ic5Rp
77FWlPSOPt8wy+eI78zHfpFzUb3LEex0Lu9DpfwVT6xZvHmmXEiom0ptGE0qnkwif6b/KQWgiO0X
tDJL/DsPO5skSGjnKtVw2O7cKuGIQSZL0C9YZVnAiTEIUw/GPtX1Td7RK31rnNq00MCeOMWdkKA4
7UTc7MaJZOTu1LW846mGqIXkdDTAxA11YWutl/L7HZE+2awXrRVIVSQ7Xlp0DIzx8KQZW9uh6bh+
mMzT/DRersvq8UoAaFgMyUWoBivgogohhTYa+P54pim2T85ABagqSNi6EuhgyXTSLBIhy8yvP8Om
Rm8aawz+ln2qwRhip8eqS2o6fXrebPbiSpiMaT5aVNbX6zjT+QZlEeBLzttH2sJDa/HerHC+zNeH
XHxXnrSJgik6603p9qx6nD/5DyW7ZQV8PuvDDn8Bd2EyVh1bf9XdgqZoOGF40wg1MCmrS/qQ/zU9
wfEstlnc2qLUZSU5ItgVQhNImEseeStAhHYJyasU4OKkDm5sbA46pJzDM3Jog8/wkHMsxksNiqQK
lP7lSOmmbTbSSNrNJ19FFrHJbIsk9p6gDQRyXpYeF6iM/oGoG7dEeAimGeMLteT+2IkeA95v5y6I
5A0VFP+vDCL6cke90cXN00FN2cL6m6ANhVHvlyJxpFf9gr8+IdkodXYoztVZ62q0baTpAnuqUDI/
VyM7D/xf3fQgC8LRJI7AdgEiJnm5EInahsWM9MUQiB0CyyuagPYXSjaf1QftlQbDGBhAw4QZHVks
/MAuXgEIBR0JLtBYGHbkI8hdRMbCr7HH5zLASSsZo0BTbDz4LjSUcK8ITOPOBamM6q42PByVKUSp
WGbQSS54llQ5inpsDq1kEV8Bv5vcjdqKkeRNe+bqOghUXcL9QmJd7RQMHwFqY34by1w4V/+mGWVI
EVQ/8DvrYIqkput4hV5sZ6WUCwrLlr3xxpTe+2smTML02IcqkOb8cyD2nizGIkGnDzOsR1S4Tz6g
VwCYsBYM6/3vzMAQJREHugpk8fXTzvM0RtHuICgldR7Sz9/DDOO5T9n1Fjiyv11CK+vTcgHf5T4z
vGSebW9kKXIsH/wkCRLgejagP4rr7vDL/qBfyjVRnKMvIZza4iXSP/i0qLMCDT5D61LzxITMITpB
s3cpS/uv5qUnZChVChy0uWlkvbykPHS0uAyotrqRbbyLcPyIjVncQuxDjwPkE+F2DekBfHRNKVhp
/s14zlRDRjfMle10qCJ6M4tbWistN8ITXOI5kVTD2E+pURQsWHGNUB2nB3U42xUr61+lPVMM9tTt
6SeZWApkM00m2cULOGGPx4YMBJ/iEeh0Gnz1sNwxEzOk+rrbUb6PqocZ/1xjZtq2Hm7EV25L5CKM
rQNsC57trjhXGuLr3/YTMxJ9vlEkPRAZldbSYLv74qztoJ37AhLv9pFUSIPeFhaiBRcdQSvrbSUk
/APwhcgk55xdYqEIIEoIu0e4eEoV22sSTijkwcQ+B7JUwn3J8v+tH/bJPFU1JmKNWUL3H73nXVHy
AFEQbD/aAlVQNEUU7wbNf2/9poLoM+dX2EFvmeN6nGjnVDt2NSUoaMF8UOFXdR5OcEMIK7SSWRBI
kfHBXvHGtQ7Ru422RxO74CGzdJVr+hunFwIeL4pg5Wm1GbMV1lqiaRZps10jP1ZIZl8NsK8lINOe
kEeNDsvJDtAwpP+jeAeTgR6MwA1PluXePoibhFbBh4jUKpcKa0ySha7F0ExV9lnQ9Xkhgrnj0Lbh
jxmMf3PA2bgDK8IDnU+UwOZdeD/HXadjWooIbW6ftB9hJ360HwGViIM7rtIJkHGY5eub1GaJX/FT
RkVUq/SDL73rAyyLoGZyWtnt1rmiYizM3KfYKXu6Gb2k7Di3r21MRvDNC6aPGqOOq4Wu9CCvAHS3
e55SjHHm/4AGaMV8e0h0NTxFXSNHkWS1v74gLzOR/CGth0s9BvZTj4wkrEzX1EF5E+5MilBulMKV
HGHxIrPB1n4yg8g8PtNLhHtIjg/0ZCTpYmkvbDVhvZoT8zBIy+dr+2wkIgcoFh0lsFBHHRoS7S0j
jmkdu0OMh38BFgL7kxrXipeVk/gTyp8jfIF3iPgDM/DlX1JZHXL42c73Y5u1bNvvEeR2hNnwXsCX
M5YFpaPFS6hpxpto1R6l4WM7vUM2KSNVH7e51jFkyMFRcOW7dbcduWvR4tJrZ58IxRhWqwb4kVYY
j4Ak2B8KCvs1Bqt2M7RhECOATePF/Y7YWnbom5ZED3jLH+U+ZgEQGHcsVHyReNN8qUjuwmASorRR
/HkkuDGX34TaphN15AMWkuHYpwgjdF9fhsLq+YKHSW2mE73jLCxPt1Z+V+I7RSK6SVAbEy95NVoD
YZTeeUrVX8dVGDrtcP+QdHmls78SRlyYkA1PRnJ4JXLeHGXAgoKug6YC9KljLJcCd1kOplUZeW+w
HNb78+bCwr2Q/t58WOru5nD+JSeqcEucblJDyFHOSCmx0E0qBc/X4/5pb52nzfvuFqs98mr/X8c2
eJzTdko/bx7cX4vmTOIa6nmhYj5xehM58TqkOmsLGLuBRJOtvFQjTPgOdC8uEnmH4G8CQapQelLL
NKuxdPG4js9SJ1DmYb3ykh2KOfhS0G3ZRNKjBR8E/g4+GvcOstORxtiaUle1xUyXpBsaHNHtSPes
oCYzyDvWhVdQG0vmm9gLWHCFUJW2E0NP22wb4dX5roRlGdk1L6PRNJA4BORXZckiE3NPmfFbZllg
TqST6HeUjAoBFKPg8NQcy7BZj+6orhTjDprSwIM1Hav2AZIt/84beScS84i8CSeKnuOjcuYWtQ2q
0ZW1wZBaTvvsg/G1j4ppiQxtQB/hNH0EViuIkRbc7FWJkUGB2g3FoW3BDpL0iadFHIT16BbtYM5w
qQGt248bUxl2/9MxVnZJzGmOko2CN2GkLdlDmD9DX57qhidE1QaPIljWf0MK9kEebPkVpF2T3czD
1jPa+9nn6qAEuJgR7DnRtNDuiD7nXhKhLFzxFu4lSoREu8MXtKh1cGM+P/ZfcSYbmEX+VZuLYM8N
fNiMmZa9SlLyPulocWoTY6YTwW7DH5L7zITp3S/DFHZgm6cVAuvxBqWbYohxCemgLLskxFH7/dvO
j4pldEjLUs1dOBuCdQ/dc98Q4iyrbYmsxTDvaQyiFV6YLqunQ2vmx9Ar+9lTDmOiWz+TfIw2tx1h
bNjMmgTDip5/xqTPnDWTs2YjiOWTELDuP1R8AQ2xf9a911YLuAtZVKLT98j75Cz/yom4L58ubQMU
22v/0z5TtSTI+Mb2iB/ZHnlYKocDXXO+g9iNDxSyJzbl8pXllK7iUtJMHF5arB7yJLXOYUQcoH+q
PFZsGZ6od8ciChWmeP6gSLbxG2LNE7UDhUmnVQBGELwgNmqqgu/airHGA+aLmuTGbMLTlaUuQKZ8
eb8h2yivXZ+702aQWllce7Om3ccf93xI27wnToL14fVgB9CQeDvPh+VyrjSNE//0sKIlbnl4wXt2
QiFiJvkYFyIL7I98sGD75wpJkTX+PoL1eHiVDiQHgn+TK8ec8qrFLIs101KMzQ2JcVC8HDzM8sh5
O3WjrlxFihwNMg/ZcGKF4ubdVeM94ZJFVl7KA0mm4X5CV85UWvruZnRktmKBiK9aXcqoucx0hkuH
6TQEip+/XbReRL6YuLm1KCPl4duoIAC3GyKmqd2MgOW5twot3kGDu9cczt+HpIiPC1K0AVFGclx5
0PL5wRWSHipBtkH1GgMZOwiHCiQTb/8cckVrkhcDSiJlolnIXnb/8cKTlPGcjRhDdM8/kr4P+n0t
QpdjaWd48TVcsHmewO4dXzN09lVV22//5AXTv51w+QhXH5eMDPbAMhE5Ig0kTrz0yPVNPJ7LzkyK
pvtYfQ3KJQQKolcYvSr+P1ACDXRR23A1TbX5GQBpetPXBehghWrkqSeLDlF0FDq1SfE8QRmjzi9t
34DV4kgFLqVhZ5R+arOx6XqVmguzvtk0nuys6Zt0mpTjku5wlPDuwAyhJ9Kjq27pO4nN6f7tWwVQ
4seHPL4yy5IQzTAKccMiH5OgRG5w/+NG8dXVByc/YcGHK2qW9NYjyn7ukTBOPQLzxBDqZILb1zg5
+n+P4GWSTMN/mYdQMm4BmrimgggNIQ8aj/fPOKC27MpGDej6SNh6DIrbW3qqZhgYWGMBEDfWwUie
8LgLOPv9W1oeTJMzKXpXxn2OacSrfCWIDIv1AV3reJ1GF5OaYLXNem1azhS4w3VNqB5w+Zye39Ei
fcnvrmNgQOTVMUpXGWOIlycRCmopUsgUHkgz6hgRjYHiiheD2dKi8kznKa0Z4Bqe/5d6XPG7UF0a
G0l/5K8vIKu5r+eWjr64+kVnBHZOYsore2Td6MVP8uvMSQ5X4VvIUmHUiqRN2U3FrM4W9OuPdKly
YNXQBgUMMku7hzDFt6VVoy0QUWBQX+5nJx7D76XhS2M7WpDTZgEBqpwUhxg1UopnwD6rRYfHPUN4
3mCD79TxJe4mKV7qzKSwNZDdTTlYzU+ANH1OTdJ7P8qgwT6+OQXW4wGZ7z8YepvbtbfDxD3kyfAv
YptbYc14tXfGNaMFyMGAb2nHfcWQcdXiCvDOlQsf/KnXQ3GedQr/gHCN5ET5nWITc5SENcwsnHFo
N93cP4LqVn5KPaJW0Qm7YRlUClmmd9AQ4MrYxiGumx/hSCiRjUIRSKrW3TZ/b8pBMRG/SvOgjc0K
SGMIA78wvrPHTF11sOrfs/CryjbjDRKwJ4+A5cOlMf26HU7nQcPvmthBw3uRTqCqz7zU2njQ3sGA
EnHjRmWstsRpXYVlHenJAEwimS4Q4uA9kxi3e1o59smzRR9w07yqmZd46Agqs7AkicfHRFhu35OR
ilxfGwrQKsiU5sKQtPbJPCui5abmpDgLg3TUIO5ao5P+zeMQ5J8ewd2nB2+slIXek/ek3EvXjSbj
WjzAPZph29nu348jkkK6whWqr5tKqoLrjeMzWexVnxbd56t4Uccefw925iSZLHN9+UxwC9KVgWuq
VQKjfWjlONvpzsgDFHNU7e9cHeAv1f2ltLSjCdif2Db5a6f7AWYTDUqhk3Efl6XgtDsiP4q4HQBx
BaHGAwRfchoYG9gb4tUY7AbuXl51P9Tbnp+95pLwLY5ADSpzG1h2l7PsQ47EnYo3uK1tqTJ69P3V
mqS/yN04/Ik2v2car9RHoUfDQ5YlbCAcjHbcVa+51ciS6xZteVWWr6SWYna1et8HR1hKdP0heA6k
lysNyYx/zU9oL3WGL2cPU0jJeL6LJAnWYZEB/zSWNRavbbSoFhdi4Uyyp1Sv2ddDFeXizPabpgiQ
kkJxsl2w00PQ1ZfwW7HaCP39aLNCmbKeuWZkBFv/4qZB/iJUZe5IDvo8SvY3W0d+2ba4rL6kWJxm
7PnZZUdkk/5ClljHjM8+tNete04FIByOmG59+n1SJsezVr7KtaFc7AxNzH4sg3ZSjRbRnYL9aSa7
cMhH/B8TMKa0meErOjfSlvEJn/giPPEt9HGOtcde5IsOvBKSQdcsfZcwayD7q/pzzYaCXtaB2+Xy
ZPlp3YmOPj9CuYN2UvKSuOU7E1Upp1XBiViinqE9IwsMk42eZLZJIoITSiyel/uEXweeeih/3pfc
vLGBvabtTiko2/Mcm2j5oK4EaOxvEwljofryueLVqDzTSbApXipvOjIxpenSuRbOi/plsUB4sUzo
bGgXBcBVJ64x6gtMka+w+xgfJ5Ms/+cdKQbbuSVFuwHV1nXwU5BJG7zGW/xt8CUlNsDcpc40NIHG
BO3HmMkbsLAFrQRp2OQBszh2hz33tyYthvh4Uy3JBv78pDBPf40yMgvYvUqbCNuB0YU1Zfxpnucv
Ua9s7dxrv6iS/THhtXXrM6FbDCQH43C91cmmxGJh0+02fG9t8JBVY24OkeMNkStsAWHDqyB2y6gH
0pUuBen439dpnFA/P4s/9Fp44onQ/uv9qDfww0SEhvLFEYbKwYMiv1YSQ5EdyDgjngaLvtMRYAPL
ACGszkcoCQjpzG0rKgxlbGCWAsvzuUppHUqi50147kdiIz1S6C0dmZcjY4V7FtB6RKdKqaAVFKrU
n2yrRUuPaAx6WGPkuaVZWwJZwHM4/IpLzsCfJO/FByAnaJiz6PQLgZNJXFOQjL+sjb529sAifEC2
MewRZGOz86Caz+ZHBT89y8Tiq0cZ8TCe5f5gRh1ze0+loTzdLjPYbORRc6341vM6iyEFHVlE6gPY
wmltizSKo15xcoEB2rc0SOC2VIO2VgTJgDwZJukWEhnkzJ6ScQMiGoILtYaOn0D3RjQVCKzd6421
YaRHWBVNg098FNX2gpbbrpC6LNCTYf1BcUzU9JPYDE2Ih6xUCUzWeBRrboBcrZ14UpSHuzG/tqiy
hu0oIz7E6i2VO3/Iq7nRh9G7MDyJ/FsgLwa7O5vcwN30o/oyttNIsq5eucbqPs5kXQ8maKUEqJCS
m3naJVAZocA+8hBGd5IuVHUV80+gEqmMAGrh7HdLTdDtq1ryYNJ7hSADcCDgqjNaf5YnxUpMKapk
OP7myp1mQnCydnu2pTSbHqfSxrifSXbqT7uXRtRUmexto6gX5T4/NhzI2eUkb5+sdEyHSQ7sbFUH
VZA1lQ7FRII12FqQBTz1QBWVDzAWxsFQcsOvsGK0a/Afia35P56vgW/TWoC5xZ+IYLtW1ZcVIaAj
V7xR01g2ipWLbooLk7qPux80/Z8/Vj0MbDpqyQ0HeS+6dAtSfshYMzQlYqzI3upjovrwlhqDqAtw
512K8I3iaOFQoaYS1J0//akYzpLNDZhx+IzwZl2zUWcwpogwY/QvsvC2sIi0kjDt4JQzODFyL15W
rD87880ME4ELGyNlI/DQQd96mxqi+amgN9Qh1URT3d45Tz28c3PPAk3FMxlGTxYoYVdLAiPX/AsB
WTg1U3VDHndWwc9F/UaZp/leenCwC+sLI+XWPGMho7FKEd1M0I7B4up9lfc9uB7HqV40EpPdaIFa
Z9BZflrQJoPSH+njCXv40rLolmtcpN9R16F07wL09AAIfGnVLKpdcUZkpdkngkG8ZWpdnps2bVCj
Zf5u9y3TER+YOux8/OhHdO0a5qW5Azpkhb4dyI/cBSoBmbABicKwr9n1Tb9Oozbq5Bpp7yFaQTlr
7r3PThVm9omOqQjX3uVTwqpjksDJB9yrnVhb74Mxt8htmigX5KY+PRdiTK8Sl4f90O0m1e+9p8Rc
CGblOeniB/Oel3GJwFJphW6XRHBjTJ8HcFNGgcwXHYKULxMMeqCC5R3mNbO7JXHp4kUCXq+mmvcy
Jc1kZHCA1I8Vfjl8IW/t3ug/OFIbFgTypeGHBnteGgl9JycQ6zDY/b8TyI8XYLjry1+y9gzKpGhb
RB9Duzd97O5dOcrCjV1m9A+JkTSk8yvOKRJyDtqaEnl68G8CCDSj3zKAqJrNtokuD5+JpfL25QNi
bdd65nZHHJ6PNNjT04jIZZNiU++h6Qyq2pUY2NtYofIwF3TiQk5VMB/1JA0KtLmzw+OXC9Mdz0TU
F3rrY+GvLs1iomDqLZoSi7NRkI5MY6nalYjNnDQAzYzMqctjovWIZXTmc6N7EtOg5ehPQ1m8NPAs
hYeknFMONk/DYkrRZnDJ24HouzM/DzMnetrSD+cVlu7j2Fx1+fAZLTyGrIHfLpuQoa+5172yOxBu
qTkBeUmzv9CZPaOab5b6n7/9EE6anyxgMRHMGI8SjekRDBXOEZYPskFvdjWKy0coYG7GFedhR2no
zoOxzjbvvoebnsFBznEgkIb6Rdor8lqN0iaDiucwmQHp9GG9pWMO3D7CVtmGKYcpF3FzUu416p08
aKhpvdLVzUFJRrAabTk03fAgJq/7ANy9hCjL3fe3v5/UN67y7lPfUl8lcRZOprDY4Fa8vLDnk9mw
PLYIJddTDYLaKUaJKfKLhz2YFGayOTQFPba/l+3b58EJifOcdq+iFeZjpxsfYNItRJQAtm9N2yQm
NBuSf+cRGCO76017qpSggPxKQpkwJn+MVgtWiX6MW68V0iVPX/7k7KciNf5dFxrVyluiWoYPG2Hj
BcLe8L/F9UzU8m54Ktpd9sUnMcirLGfeRHeu28KOQoIWhL0/skTg8SAv2QnoEDrAfUiJTQnmlfMf
DB6gwqrQckN6s21Z0A/voWDrSP+ygBV9OtTonZsc87aT7pSE8ig8FR3nBxieXsWEYqrpzDQKNLsm
PfkkCDrcnvh2Xo9Gu5BoPN4OcWXIEV8XSBbUYQ1CGuzzgqBZIaG6L/Rdq9lRGuNO3laaFG/8gNH5
Y7sxbvwX7COMSm+RXk5LGWp9AM0y4OtmIpe53Pa5wYdWqkfD3NDYnCs1Lmu7VVRdgx88KSaPx5VL
xeM1b+wtxk0LIckYXbJJR1fllqWIV7m1KHuaJoZ3hCfon5PSqyK1d9re+9tzJ3h83k6tKZCmfkIl
V4GD/7rL2sSNFlOWNRYEr9ahMlP9lnPsT89ybvND4I3BTHl2nh6V5JEd2MitxevkCZGr4tBRulNA
ltx57mkrYlVBWw0iKoJu9EFMY4rZ/vsVv4piOtyXQGsRx48GED3Tj3PGrgJWN6VU845oq0E0oAYD
XvAOuAezQIBdPaOegIQR8TR5+2Rigcajbbx0bU/mvb7a7TU4qcjfQmSQxN/vBvgjCxQoUPGUkJTd
50YPMPEhy5zWynfo4BnJaj4zBGibN7FYNgYXrBRh/Gzu4v1sKAwJ369CGxFQlRTcY8LK8XyHKEbA
m7ZokceYIMvI3T4OSdHqEDRcOwwAtasS0q9Qmxed+wf32V3sGQJgTx1TV3GDCGgyCLuixDId8MwC
NH8Jr1vZvchPH1FL7jEWDZBmr0GBjTXW9l0Xp8S6eLla2hCOAQ8GYN8Z8+W94xX3h+Nq4b0XTqfT
ySsIMxyj9HrWgYIfE5SUzjzX3PCl8ubtE5zH4NJx5/2iyYRPuct6LBz1o6oYGMrcYfuT/n+ylVh7
ckDdk9QHsdrXrsI1wsP4FpmDLsWKALVDf3D0HhrydFjWu3Bv3yheJTlcwVik0/hsHeKUQTY1kvCt
17Ryl9lS0FiT2u5bwSbScSXc2orUTe3oETNw99wyaslKeVwHc9mF8RcNQ2EwWZo4g1xAbfqpz+Wh
D83haVS+6LbNULMODvOfUpRxDsWLkGwrAtFNjbVkY6BW9/V37fQLpbaTF4Jl1CvsndbaLK/IYH8T
XhUl6DCS1ehPnA8slPwHqGs+MCh8aUKiFGOmW6NQQdCEhWaa5MEwZqg4el4bzu3FqNmVCTLPeJnq
D8g2bxEzYLar/X3Hw79XFdJgYQdu3DLFAvc84JqMfDjezQo5A2QlsOOj5qMPmjdg/8wQHmRdZZfZ
trlk0mfg50dvSk+Ezp1cR+5+0ykqVmrm6EEWh5USP7K0E94wOykbc4gRQ0bkc8pYnoElbk2e9v2D
GTIJvfUou1CS/JRBe0Z6RQJsHSrgSeOmvIDrcFS+5wAIXRScM4VqVHA+OqEyRWPwkd1RPeiLzIHp
7w6d9UI6OCy0/8lNKKpyDniWNuFOiFAQBjZrf/W/Ww69ifJ0XMzm36hqksk662Tik4WJlR+zFXGX
N7o42rusqvso20iZMmDljyN40vutbWwpq40CSKgGBYIjgVuAeQA+ef7ccjcYlPCwyKZ4CWjLDf/o
eVG9H8iGd274M9x4/16l+IFqj6nBdTIP4vP4XDSVm8JL6K6fr1k0Xqfv6Gx2IQUxJa+bdTpi8eIZ
I3NgeztY4RGyMWj08Px/d5Zgh5WE2f9ERc9ZnsZulZ5c+vYZLWbuetW7bTWDSZSSgT9Bdl4RnUUh
buBH9QMETiEYFdAqwSSL/RNtaARj/VONTBjV92JyF9DBYdMx+DtfMm9y0DuQaxWcpkFW3fp26vZl
bAeQMcrxBlxH2jHDO/xa/fuaR++p0gaXzG6mdZ/F6oj9vQhcd8wkNdTGUUUmuW9pff824Ttc/D7r
PTkPqsM33vNvky43v5OMA71yYIQrHQ5DM2O7D2CB7kElbwY3aFeh4XnBaAWsPyZQ8KnqdD2o43zj
5I6uZfDwtwW3T4/Q2YhEciECihjjdPH2ZjdJB9iF4BBS2mvCB2oYacA2fyK8sTtCVSYzyixLqTXa
QhfayKpzv2V5ADy7b6tNv3vCdBSPCO2VLXKT/AIwZVqy65/6oXhnJftGXEQSvsZj5ZbO/JKsUhfh
B3dakeZt+q3Mm2xIMhJiWeqI5XMHNUD6BVgdmAb7BKaHhKuDOZhG6hosGLm5HDoRHqDgKqaT7aJg
lvFrJLx1gkjZipzTnYpZwlDPLpfJRNppI1/jn0RP+ZquVhjsc5gvkXiUaSk+sefnp7ab/dq7pQhy
O4IZG8yVbiNPkopoRKlXx3v4UiERWbzatNZmh8MFCUZfEK3ewj5VQz77C5kvcVMhIjNMs27Jrt3v
LbvMiY5wfT6jM2r+fSU5ckCDXJbGBV2IwVA5J495Cq4u7QZFObhavqnDEXqtWUw8q7FpiUO7Z+t5
YFzIUF9cMbrPWdjA8Gsdmk0RAEPUrILDd6kW/2MyMcYwrv94ntfUr8t5jlMNGix5UjKxL7E6r0iA
aGFImiAOLKK6zYVmnNiUuvlJhTcMjAY3pFvC6bRmA9YljrzoC8TXKqFa/bGsfVfpNBEIT2Q57hmL
3GK7HQjk3zU1Id4AxTfmiBjfEFRDf2qwMVcQvA1ARiG/LT9FHCKbF9S6E/83ShxHQ9cjnCZ4DMrg
eBu1brM6AaRE++JkBPzKsWmMAwan8da+wzLdCbs0pqmrbFJSR4xMmZvRi2beflVHB6hJE1Nx8VMH
Xrt1S4jSAIhASRVTq+Kt8c5nPAXS1ypyaQaKvvGYQcw+80QRSKLFqGHDu3yv4DRJLMCnoN50kdf6
InlzHNyWO3hPvr2gzhLxRY2MM4nRzrIwCNo2947SRnRiuMFLryZgzSeCaS0tLeCHJSd9VqKDHZ9E
Rh05hqEGVMrXgCYgO/pYoS0JeSohI4xlDDs1N5zNglLGhm87XipFXumrXNeGdZXndvovkwnXM48F
RmxYdJWlhdKi9nurpVQSPBpBG0GMRi5mse9zbuj/+d8Tao7rcNBxofvekUT4drmONHqor5XZA87A
Bn4r2k9NUmDwCqTzdMxRhcwturQCinQHu+lIe/oI2zikyORv6u/K//noZ4DwSrubdP8L71/QXebn
JIaAWHxFPIb4VET6tSpo2Y3gv4hk2xivmkSTRCzLUWL97CjRjSMFDTuwX/kdGpZgWoC0z6qEmiIJ
GHfnSNm0oBkN0Nn1wYyo9EF6ctJDIOTJjW2qySdop05H3wc0PXb2e6nJpmYJXBzffy7RuiBDXtOy
LF+lAmxHATv2BkFN42HEslhnT6V4ljy3hl1E0WsrK1QlxVBe+jyCerkT5wVQpqkNEwg9/+e+HX48
e/of3tg7OsZru6JYTutZ9qyFcs6WDjHWfRyKmgnMnCnHbT9IZj1cwqOHK6tMaGgz79QoU5P2e8Ut
D8x/7IUuTQbGT4lpn/fosb0DyRxtNXgIBnZSBihnQ+d4Z6Ox2Av/6B30gjbDwH7wPXj0EdD/YQAv
xxJriYst/TYYR1bsDjdM2j0jtsO4VFMhozX1fIk/DJV1Xa9k/e6ZBPZoP/HAKfGaUwj3bjrHKrGE
Kxn5Qjet/ii2aL2uTVe4roN+vQRpEPm4D7X0Y5tcuZNEXDdDM87aCX6AHpgkAPmoyMfW4u1KuTjJ
X3YY4Pf9Dw8KZlbCbHpLa5OGb8E9FzTzwfL7dWyjZbzx803eOo8tw/0h4T2At5k7mnReA8r3Tp+q
8QR8OrRArhSXmRXDdly87cU7TtpjBt2wLh4EAVsbD3lF+QiBqWamtEMtMo9O4Isp7uKvO/jSdWE6
HPZR6tR7QUpWT7HA6VXYqai5aFK3NhhXjTkMQZkPTNMg2VewSAQJ3dntLCXtDc0BHN3PP67unSFD
NNF87iqob0pCfaANDOIelY595z5Z6RCOb6tEBszhXX80Kxyc/V40hDKUhJ/+f+2HBPoXaac1zXm1
bjvwI2F+q5SKX6Dxt4/wPXfji6wkj9lCXircVpq58F0A0U5o9kC7iy0CySU9UINsx6gLAdlTD2dm
9g9aRTdrJ45QJ8pwolM295YWroZBoOLRoko2i2L83EVeN4xENWvDb/W5zp0y78rlrZ2MRp4vRDP6
gV1E49aQgqco6tbApr0yDYzggUsC89UqSCZS67a1mv0t0Ewzrrp5uCf0+Ln5OxKxErKSacXhsn7j
/NUIxXIRpnlbSzuUrQNi7X+0AsgPyZLM1hPEaCOfVWd3h7sPxau67gQnCUirT9G1ztsIDrPbSRht
tL7EjHCR+vhpyQcRbgMv96qhrruqKKmICbO7tY6blP1TmoHWmiIP8TVdCnYdOGrPY63fx27UazUk
5CSVrSsN87fExMgFoD/XuGAc/7kUiSmoBG4Y03xyCWgKGKFExbMD4nCZ3mu+6MM3tz4Q/2WN8/Uj
rttCOCHu7UXT8v3vS/5v4e/1J9aKB83OngFwhEJdOsIYAyfAeU3vRy6Em5sUQcOE2fAs6ZwiYCah
QxhAKaJIfUTK8Z6AuYX3sjZ6L1T2PI+NgTOWScz2r2ltAI+Qogq+HSewqRY5xLIn30H+J4/29hjh
04R808l86nx84jMFM+MkbTtOFK8vqzSE7stJ5EM0IoadBu4n6j7mnqLW1ifnldajmP8wjJ4KQo0D
H2OFHo8KFDWyOVeCgoYAbBneaXePhImJWntran6XYRHOWrtYpRTURBLpHwulxjGDbxnUu4NIZEbQ
TwFPxQZhgTqWiHaOZyNOI28NqfE9IBkdrdpmQkrk5DHsqYp1TLQkIfuJi7fyOJ7tLUhqXwlTOw/h
Wd3cdTIYGGyXRFwe3PAmo1IP5Yj1b4sTXxQ7Qo46tMk6PiXDobHXy6QDimaEk1/JZ4oegEtfdHC2
vaYlVPVSyvzZpLQNp7+hAzE7DcWM7PiZRUdh+wsxfhztTLDbbFV+fcXc+J8m7saI3ICoMo7LIe4c
YjJRmlqpXas/cuhK3QWlzinZg8vTSNwo8M0KNUPnlyinOzjIUJpqap7bAMvPvMK+waps0KhEXPbQ
CXExB5I/cZ+xM7F0en38mxUFe3DCR9yorK3LZ069cAZZixvzLE3zcDCrcpNMc/zRmDNcU3TOE1zX
JSW+oTQleZGYcHAI9XPOQCKbPnM4WyGeFkjkfoDbl90kQnqvCuAHg64ceL+EsLUbb0qCFppENaU6
2P3C8tDvQWGuDPcpm5GNu89n1hPfIaHaLS0rp/khqQ21VbCnKMl8W4++77CPKd/ZT8gErpwYX4l2
1I6gLfDJBPtpBV0So/Xu64EbuskqDdGscgb9Y/1BADcj/udynPoBr838fPRYAeQ+X9aJxL9OAJPU
lff1CGRdefVnjzEynYwUmofGh+M2XGJuU6h4sf5DrL8CQaEV8gHfrDWIGkUpzFfkysiVbdx2vRzu
/of3fAY53v7f7SSRsE7GrwkIeqNOUyeUwyy0Oivehz9VTA2DLMg3+WnVG7XqxzpAFXnH6RUKR3pP
Klv1f9ZPeMe1RdaUGNk8j63v7MVbyNJ4Wit3W9MXy3PdobROb/7hJgkcAOkscPLUO+kTO7BM9/mN
CPBQOicJ3DKfJMi2niLwgJ8TYfuL6bfAALAn5cWtfrJiJJ3qkmAlBtxt4INhGqFena942VpmaQBX
2rZ6JnoXQcwhxzw5N4KEm4rSeSU6szLOEhep5Fk+IYIaXdc1GgEE4iC/bLEEPMuipy0TkertVd+P
YOb6vkkk515MhKZ7osPB5Ep7rnf+qHyj2lOGqO3Bt+ii7AKplKpcIL8Tw5fiMG8Y76qS2+4ug7n/
r452Hk2Lp6JX6XrxDUkW/q5yHbEgqLBG40VE2gUaC6Cumj+WlVE/LmSVdfX72x1D5/zN/qlsJN66
XWquEJkc2bJTxJy5SDeyCDLjFT6np0NIyk+VdqhUgDxz66HTW1hJJPswGln8zX4UMdL9h+fZQzM0
lhbte82NIdtJbVFh/5w3Gsl9vLxO+HnCcg6wBCP+8ZXNU84UqrPeKylmgZC88we5J6LYmGLuT/2W
sX8qtckJewZ/hugQyua41v+yOywxzdD4qHKTBa+qfEUR7h8KgF06JUvp212DiXez7DlJ8ePV5+Ex
XSQ6ozIHFNTqLo/wBMUKip2z6BaUoxFztOducMvePRxc+371j7U85VZJ0LyT/+1L4elAktOIMMT2
tw/FSCwQrkuQeDSEOi8qayViEcguv9cIH9wWx52avccrgB897weOovLWkw+NHt2mbn3k+3bU9JZW
MFa/Wp6iiIg0WiedSDNSuFuAbR7jQQ5LDXPPfXeDb9z1vu37e6MAvndQ2SaQpTeFtxeOxEAf8p6X
R9n/bFTHogoStfGR42DKtPVRkY+4GVoWblnEaBPP2nFCSnnRGHmMlYqnGL8M6x0elnWSGXg8uBmr
1p1FiWLa3VQQlxfb6m7JHFhOnlOXkdK/ryUT5fdkEtUKN5u/GHdLxF+y5QBdqv6J4foQXlZ+3X6p
7FwQ9am46/8i1OyOt6e0cgjNmX/zyLGlEF56/Al2vgY+4dS/pXlsOMa3ytxiGrkjqYBKtYfU7CRg
gGZHV5FQJxTDdOV/qXZ5jnjnsvg5AHk4XkXw9Qwko9QSXF/x5sSxM5UlXHwALb5y9limLhVq8Dxt
6iPcgFToBY0i6svqZA05ie1ItmOxirFbHtWfDDhLusIZgoPtUTcPqEaF0dEIY/OZoqx+D8CGrIXN
8uQbW+d8v05vbCdkBcE5wRqUE8P/qNBQoCd1RMVDagNBE0Dskwk0zq3EiOeKpWAXHoio/gSwZwIb
afrxmwWEutNF0AugGBtnCArrDo08/8OABg6LJIKNZKMyELG8hFb5vk7qE4DoHmQe0hpwq+0OKt62
cdDR36bWbvksL74S7/3fZ8vCw89tCuOKEckuT4ncZDmUZiEoqTJNz/NTU2Fm/wMumTnMBlbHd5M8
ro75KBMzyCaqKLCQm538n6ZiCUmHIQrOcQWIqQ9gyf/EgvaYOJXNdOF2m4ItxYA8WkL364AXVDoj
3hVY0ksTZPI3VJLpCxg0EBEtXMkXbYybRMJ4+vl7+xL1V1xHT+o9CJOFV+VPG0zozlWI6n8b0nIX
P06giYMi99NXfn3l1tWlSU+zt26NnkZ3ymKUouMpQU6w66fQMFm2zOSK7oBHMOyW40qbkrxk5VO/
TittELQ1dNZi7ovjHvDVKMM4Mc+ONZWdOvZCCAa3QM2JT2JxVurQT7raUxQvA3JXsazM+18OhcOE
iNFcCn2XlS7JEpA7W0Jfb6qepZoYgkI0lfpTfMiiwAN1sms2eeSaCqq2G5cav0KHxM/qjk5G21Pt
J1Uwb6DjSFZO9DeM8nbbS/vdlZSjK4GC0ps+TlnYqgFDi1Ky/oT4OZHsZ9W0Cp9hNcd2RAz9n6z3
oPTXNY/5gFdy51qgJ6GvasY9GUDaiYIhgWG8Ov3GT4TlOLXqBYs2MvRAimJiaMqUrm3cKeRHUtTV
NyyPMGUD+zZZSmUiYbTKNJ0PahG9kxP5lD0RTbjFcRofwXM28nPkJ6THYKPaLQTt+NKXz6JLpeVz
GjvZnKc7K+TNM1r0/pS6gJh5PPaDWp7uQGamQxw5i1MBc7T0vIwNVIDzYdsNzpdv/tDroxGRSuV/
Db4jKucaUn76FAkD9dA2gjmarIyF7UtWO8QaHcurJ9G1ahrUDBt2pYHvBbgoX0CPoUOtTWGpJmkV
Mcx+2gxuJFjztd6A2MsYW9SC5bHj0iEp1GHsRVd1XQS8w6j55nUpv2XO5/UoTgJbv30b256jJkma
QpucORLfXB1hHfu1rXyKuGHNtZXI9cFlpSwgKJCpExDaubKQBCz1Rr+Ez9LN4d0P48jnabandQbj
OIbg7lq+nexeyIUUWF0MYq/+0iRe9j/7yWaDtzFi4iezVwQOjvi8a5aL2WZK38XtZvqGXKSSR0ya
kgzUiIwbYivqHoV9xZALObpHcz19NM8C/ldgzV+7vmiJXmL5ZcivpR50iXK4k7LVouMwdq9ON+NJ
1fhqSmiyO9WsEU23LghwTzEU5Bktlet4JZR1b4BEauK6XbzNjUqagzzdqkfim5MEw+q+Nh2NTYRd
u+RPQlEJp7DT+tco8cPgr+fTCOD2c7yu7i8mJgYSR4CDHx1+XsqlhdiGnxAgv023+QhyHdpU3jAq
8sPvzvinw3E8PHWSt7dB1eBf80ol40zT7cIMDzDUTnUWagOySmbhcxIExtBqZRlc7hs1+O7AEWhI
WyVsoVQW+mTvnDCtd7kXwJWaEcNpGk/K0azc00u1rr/V+6KAWNzX34Fl8Yue21i71iO8WUzMCeBJ
Ezqaqj66z8tFu0+zDPiSAv9zFvEBBNFP3Xslwnx5A8q8yhQDEY7Dk7ZRfYD0HDABpOfy7i2dwwGc
UvB3UemOhP9p2b3msabuqE6ezFYtRYir6f1/kmlZaQbC28ED0cXkKQbi7L5ILatrBctcDZxfDljj
vsPWEM/t2O3M+KJZ6Idzq9HBkj8NLyckjbsN1CDAg6W6GVv2Bo6Sg+Q6k42JjKVJNbabqag5CzjK
Az1Oeeslr48X6odvAs7PFXddtuNbv3BXrpoYm6Sg/I7V88PiMUktnTgTTJlNKuBXtkH0pP8aNpqV
JQw2DaqNy6o55fUwcyXjbLVeVofAaOjU+Trci2iq8dZkYuj/ozrX5XHUdopkR1rrUTSe5osSa7bk
r28fns43IHXRUmUG67IPPwjRFHUvFV9loZLpQ7+DpZL5geniG/DseIHsmwiae/CKddFfFyNvpQ1b
SVKM6uli+SMCnuPEc2+YYkUCg1JfmsheRFx77e+sQuYAt9LAw/7nptNWwLK9AcFkUE2pGfEQa5O+
BPm+Za1kIxEXNav/XgJ5tDRiQc9xF9xMjQqRzlm5Mg6AdnNeLHX1RpLhr/GTrdgkDZKDZVHjUBXh
CtzJvyJUVRMKCy6SLi8MGmwo9ZqZNtGum12d9wZce+Phv9Qku8Ja+3yUw+rPdlmjJtpcU2zjTr02
TbayNhBzwQRkblHzgXVHpwSEr+IPW6xoYoNHsZijSTQQ4tcjIRX90HA7AUOEqdodlmyiClfjR7Iq
Dy47/LNhVvXlxpFSD/C4GBEq+TJdpnNMxWB83/MP2o5Rs3cNgCiKYHc+pkvsx8bfeqVe9Ar6PqtL
FcTHJUIxHP8QIWFm2qQtakXHCxGxHrbifE+g69TFzkPX7k2ZOqSl8RrvemYX7E3JlJVKO+mrfXXq
NT/Q2gtiN1R5lPtGudWwEYgi7GV47sqdXe7mNR/oNJOPhyHp4H/QZ9VyZFNsdj9aLOR2T4bTSHyx
kOg8CigTfhZkQIzhjdMz878m6gGkKOADrdLaudyt4Q0OjpSIhodVSVFMTAsZv/TrC8AFhT4bJjSE
bz7y+LdbqoRAOW0kzHGRwdlZIko61e2sC8EBJqsu3RtXkfzn7Z6PUgHAdzpX9MvOVd6DfIfvPAj3
zVfhZxppWxCRLHFdqYKuKtPCOeIycvE1m4x3xsLbUlDJq9Jaqo4yKx1E8v/uWZRXXPiNWet8CMMc
11FSgN3/8KNTtR1jUMU07hURG25aipaFwVzypxs7BcSp/4vvBPwRkxWxD1wT2/7Vo+D33iWz48Qt
hN3STwodbiSN3HB20BIstOdvDI08EdiDrH/RUGDMkowdtjOxWNRZtORUtFfjQKiBqJnraJo5w9zy
Hg+0QXrpPBm3aYgKmi71J9FPomWaE3MMhuwo/xu+tJTuwglEfgo72dHO9vbEfQkDnIWW/Sdat9IM
GR49D0hiSCBQkhN5gx4s4ppk1yUn2J7F4pfePWYYaFFK1SF1LK2qbXs8re1j+iG+ZEYADCHldd3y
8hkDRLzFzu3oHYDtGZYR7tz8c2JvzMiM9XrMByjYVpWR8u/4k+7CZDQ4F0DWpQGmUuFTkPtMrnij
v/8DP53YhHcxnvozbfk63R3FHCQmwYjeRAEhj+nEcZBXsP2kN4x/gYBvL8AinKYTlUFbob9tKSZ5
z2YconxNQziZAPidsBcLLdbip/sR4LEYU9I6pl86hLKLGa7KmSTiMx8XC9xDzjLn53+S43dZ1HWz
/B8AQ43Kfs2wfBan77BYeB7RCbKamXlKEhJfjfjrHbealY9eDLQAcKEGBXQzF77JGqS57BE2DzS1
8jHdS/SbqU+9x8dBUV/qn9wtuPojyv6pzE0ggqq/tMkUFi1qJKTd2xKFE38PbtEVReuA/60cw0C3
rKB1C6IL+UGABkx1c+c0yUGiaoqO0DTJ4fJNBl0ScCnK6dXct4qX4TDn2qnUkt+RpH8A7HU+/IV5
qvJRPGFLdQKinsZVs/h9732T0xDYFTLLHpZgQ7LA9AagfEvgNVCrojynK90ptU0oHDDYWA3uHTHZ
JK8W8EZQtemnvbiNH5XhLTfUa3F/KLBmX9F/3wXUIsbbHpD6aAfWd2+XAxPZc4pPjMRYs5K6DHX9
qnRx1+h79O0L33qaOWVs2ihKLfZRz4CtsSZQ9ya2GxFFAq4vUbmntLcQwPeHAg2Fgvm3VZjTLCkV
zyLyNER1yjzyKDnvOw9BgpJIi7QgpS86NgLghHvnPN6BiFUrQW1XwG9fSS2tgdqQfojr9DqOUBsg
8Q9UJ8PZ/wMhRRNGfjf+fR+AZdwInGjS+NMBwHSb30POV0bGxJpnraYopMKIen1IMtuqkHPRTB6O
Kwlcbuzy18haZw8i5HHganZasCs2JGqmzQ0G9hfEJnk8SkBY515iYtTjVF5Kn3nmeqr59bOU/ZkJ
AysZnufu/Q8Ma1/o5+WIcUiaOW1JdVq+k0cGdFeiiqYNs53YMJKWvZA4uvbPqa3pMlQjbJ6GeTur
yfVSBG8NmyDYe2LvRQWupr3uaJoZOY8uUEO8aHDyNCL44yzO37oD+u6nelO5BRi7Q99pjKRqJWZb
o0EDqQ84RAUH8kCd7YYWvaMtIZuZiGSFXc+bb66qLizxnayqk1r7O/pJboqajnZfoo0wYlRM6eZu
044Kmr7RB+PCHotqyrT2vkQKUsgRYODf2wawiLmpuDTS38iQl3X2y/xsQ7KIRbXqI53b3lCPNBTE
6t9ycwPPAK/FB4ZHJhFAIlPbSCyApnYErFnPz1MpAfB/2EBCjU7jMYaGJJwn9RtZGEZnIczBr8y7
hblfZXDtSQ1RBk2XcxvE1yo9wsrcoXmklkp+wmm4xfNBUvGVV0Tqrq6k5t4uFyJM6OT4CEnYGH6g
tgdgeCGLmRFIKxT7JKD/tBALStDc8LSQfgcItzzQtYgx0f+EUQNmUg+Cl15/04G1PYhyC+8MyaNr
6eQw7PKUR/LnVA6EFY0jWXcgpx10q9lyNG8TJ8Js+LnRPs/Aq3yl45bKvEofZw1sT+68Qi3RFfSj
WY+zMmXVxZS8u3dFs6A/19qfhEKJ0fdq6TPazVNqK4thmRCer8nFg5by+S6BJo9KrTgwWJhSg7FZ
ddjVtdJVDCncX0+4OIfiihZjcXuWeUKxA7IOmA26litQZEmwRv3UrQS2sQq4s+RFUCdwsP8gR0vb
4sY87vBdfdNxIGMD3kqFAxRSRCDDioVT0dzNEr/XxUDpnZb98N0sHGIesfrL4cGO6MVR96CrWv02
VvfKI12uA28n++N+kpJH+NeL/bTW0wma4A0ecb42odXMVfNygBCM6Nt65Gj8URuR28QLuoSt2pZN
8e/sq/sMV7gXce1jNZuaLaHpkdJAJIzF9f1Cld/WM0JbGSyMbvPQ6kJqXb/E1l3y3d8YLpHMQci2
3RjIzPeLv8w9r7lSrwg6p3G21lt2AE4BjGk/iN5euz+Q5kyPDJKtvXr9hxc5edXt0uDyLVAqpTWr
CIOBzWSFPnekYGzWPaZmSL16dYu1BeJA+9dFCyYsxAWe3rUFWAEXE/TCD/FoSpr5cu/XgCtNzL2N
pHKsXJIfACKXyhQ5tSfV9GGiYWu7ti1Vw0RGCcTKI6MZE5SMXzLTgl+cXdRl3wEBZp0tvSGHDnJc
iJG0phXijYm3Eno3Lu5s5tFh+9/zhfRzUUmkyCz0SgSHjVOb2jv7MOAvF4uoLqJQRvGSszeHJtIF
YygfYzFAcJo/jdbYWC2pxzorUtgiNTMjisulEw3jhkhB8amEDSoxK9wCTidWqJkvQRG8dojxQOon
yIBHusb6SkoHO59GPm4KBUIDunYVgLb+MUEl+Vxd7PGUf7b38pxop1IwaektVXcodV4a/9ZJQpCn
woLfw2UEuyB9cajSrPMsO0AEuYG8mSRI6vwexmCcuDIROkIemwh+CPXLbGUiiCHYa37MGYx4TkWU
OrXLlxTmnCzA4O/SIzRyv6+WcFs3bz3TBeLTxSOkmsrP8j1Wo+1F6wUWNskJJdlFtaZL0nqcf2V3
ry9GA6iSOLkS+6MxNGb+TF5Xj5UdrXH4LIvJczw8pe5OSZl1+sqvRMRgf1deuI9gda1TVa0iscNI
8LA/pFG3RTQALSKZuwobiXC3nMoKaEPue1WE/yyEOTEnrkGQmLvrfXChgeUolJuIu5AsZRNFkV5A
bsHFw+XKLdP/ojf/wVKCtNK9KutlSxIv+8YYG+Nz890TrIQ11MrncehMrBk/zkmEmbqMYE2cf3J1
6Gog9GoaCbdRoqaBz6hPDlJRY4IvLUR8CIzkLhRKL0Ud7oyUGMiyW/1VfkATxc4unvs/I+ODSpJ3
JIzK26dX5KEdF9+CrtAc6NT/Kfzs9oYAfWrppRqEZjHDMRbGpTOb7j7U7mvjQpPBsG7bJxqEl21r
cF2YqpbL0eY2jeb4Cfhk2qd42zfxfg/CwovkMw7gt8GgptuIq++hn/uIOeQKm7cJwA5wpZkkedB0
BEMm3GUo3jlx08ZPsSMGRs9D9ZDekUTl7P99iWfxMUy8hcor7+ypcIrMh2dJ2I61nKAdk+gq9mMS
Zx0jdnLp2oYlBKyxL4ooyDUbnkhcHg3qnGNA5CJeq/TuZzc6rtL+uYWLY0pvSN82iS5HK+8yvpnv
Iqn+7yQSnM0FtmngDc5FW6+2K+oajL/ZQ1MLqGeBJCqL19pOjBrK7gnKq4S34IGgz/F+rjfBDF48
1rx/ylCwwBrrIPB2WDxaVKYwUzCCSGNq0N+l/DOcVR8Gtj2TFHYWBnKJX69xeMFQgqF5u3n9Xi5N
+1bDvEtUptMDn5+KuT+g9tMZCao+wNYJUeFak+mLi0jwfNT6zGzfhsITAiaqLrsnZXtJKsvc60h6
yZWoO/AIOSHvDV5Qhb9b+pQGoLg2XtHePaT49rQK6bURGiaFdxLinoZSWTFOTqmaLVWll+vsdtV+
5YvDkUvhgtcrAcWxALe3OP+2v7wV8qxWWXp2cWlOHE1zr7SihYI1UGx9nLiq+vMH4za1eR0hpB+O
MSfW9490RSf33TDD72NXugo2t4Fcv5q9pZjFdpVRvQ99mMDy1WDY7EP1U3UAyToKKEsgJxkqyWfc
Oq7+SFBNk0rb5cJBkiMRpzRHGwbk11zqueEDLsg+ym88OK3/9NLaTaMplblPXn4rfOQA8sI677y1
gDQwdih2Z05nLgdjQi68E575rfh7stXzFZa9AOkTDg3Z7IrBN1c1vCSWVT+4cBd1sAkqfu20KlMy
M9AinfJ3oFGEG165YSFBIF2N94t1QqwUCj+8UqWX7+ua+W2j/+rcC17xXaNqH8EU3U1CjlD9XMWs
1OzSOW47E90nAWrdu0kYnXHXC1N+nL/LKtgts9YFo95DlimyqXUf9imhHNq58jSlt5tdXg15ZLHB
rjHv/SfnBRbHyn/MRqGmKg/C7+KvLRFGV0+mMxlxXsy+1i5EAMNBoruToIZpx/HtdqkMM17WQf+f
h0SPxiqi/G7dHemgY78ePjKDHf5/PFzudyY2/oknlGhm3hKC9Ej02XTlX0BEExyW0T1b2hJrOfuV
MWPMMM1+1H8MbpLrcw/zDEahmZXkUGOXaoH3aScm0rkPtaDX7UgRhdZtRMwMrfoJQRFHbrdXqPQk
uqmI2qvW5PFAtJbzDr09aDk37zz9kefQmoxJCzR7cOAWZ629IEUPRtk1Q5BVsNs8lnu4jETDxOFL
jl0KTj4Kh/N8m+ulvkULSMCjqb3T1HefHIbqiAqjf9sGMgnbwY0iZp/FQDaXvxB0eu317muk1iUA
Xmo1L6Uc6bkP4nzRQvDL/O5N0AYhcsyecAPo9VvXWK4Xc0RN6kBpmz3KKQw5uIHwMbGOiPPtBc4A
4jCRKzIrc77MCMt2+vFMaH677XHV7wCyRdkRYuYYww4tT1fkaILVuAx2sCvPgaZDr6it++joCSz8
iICoESMkdYQbycqq02JQje8/wpBLy6p4xPSGXXJazaI9ROk7EbhDQ8IJctUHgYuuRJ+cCja/ZCyO
DbveXLzQ/jZIEAGTEc5kZJWMmDOWW2Nl3H09cA9mMkagwpGmf83Un3rZNlmKSVogDYi2JkEM5g1X
yOnbGnu0hcqONUk36roeSlwAZsGkQ8Ehab+J/dMo9eBEWlJ/totGenofutJTXG3ZGqWH3GpCk83G
jKxpkySI76HXbcWF/VKdWFwMst4UwDLw+wSDw1MSoV3WZmf9YYIHhkPXXdwGXh/LHvHe8nrEiFZ7
FnlTjYMtRblIrP8LrAHpVHHNp/4r71Tavv+ls0ioiiQoQ6FXvxN9ujPrVlwsITrQYcG4yX/wLv7o
6A/qxMqBzDdWp8Yqcyp5eHF/r2DvnYK2ka+Auvg+etGqjQnM4soL933z6CC6q8CkEI57fqfKMcQi
dWwys1VoKOj2sfeIX5iMIsbK0cRnig6tRc8HDGFCXEVBJgydMYd5RWUDnNiePX0CgOzm2Q9VKeeI
Sts5iYapJ445vyXFCwHGITYJSd4Y106cyUEJ5oXIYzPIGdDmKlliIISBM0P80YQY6wDMz9Vg4GMC
uV9ai+/RuauvQhGwhmXVvL/x1no5Lc3VXhE0HEL1Z/n7bpY5xoV9y00XLob2AT381MAHXLQ7w6Ud
0MZmVaGVKtvDs571N6ypJ90kqTmv6ysY9+F5GG2xChlvuRCBMI/C93IKS6kZbCMPn+GWMdAVhWqE
lvm3aD6704IlyLsg+pSn+6ZJUozGsC/7Zue0cVdFzaTZs1JZnH6NuxlwqfI/RqJeHuTGKssEIuT5
dRgKxRAGA98NI4GSAwo3Hxd5s2cRySt7BOuLAJuu5xSdlcW+nM+2meCKKsHqnuRaYTF4ZgW0GqSh
f7dogxGb83rxu5xWsyKPT/m1wZZz2xWtpxbe+ZRtU91X8VQ8MjuUyPm33Ox0XKbL5dVbHD7BkRkS
JnbyR4WLeyWGe3p2d4NQsHLI3yNSjiD3SO2NEykF/UdXexquU9yP0lzywo6o3bvZXEgWQuJ6iQcj
7vla12KERgMfNZuJs1vQti71isHIn9aSej4ZAg6E5yUsrer1XsLsT2YZkt0d7oKGjTjEw3JAvxP/
DVXPPM/LiTV1+QzWSCLpe003LeRe1oi9a4X0HgoX1bnewC3Yz+xcm1CEEQc13XbiBVPGhmrGGmsN
IPAKh9TCkaDULLCqETTXeZSg86n/ia4qZpHYOrbtWKRgqoUZbuvjJtT1yXZgN2pFWbyDykBFvjEq
rTbtRxdLyY187C2/dpuelualDjZESQ/6hG/7uVptV2NCRlCrb2JUGPj91GSO4G7C6MyiHfejAD9w
w425GWze7Zak8cb80yywRKD1bkWnmp1Q8ERIwahogXAMS1eYehJvoCB5cvoXVv2K3gdXAIJgH7j5
dWRhjts4FVw3MjGG3kKNN0hlVHNUGV8OsLR37hANUb2HOBJ7UTtgmOpsxqJo/TJ9Cs6plzzrEjnt
NtJKQgRkjm0K2x69YBqW+LiH8kJd+p00dx60R2bHNqfh/s6CpIQ8hMhvq08L6T4LPanO/muqrxxA
APUFsee/X9PXCg50XWqeog1P6V03fTKO4xGroM3tuEH5Y0G8eJApjtploLOp9aJUVWJCKVVXRQxx
vn+8b/v06TYframAOesh7fKTNg1QZJHmbPISrv6raDlUwhR7jNsWHN7PToYMAIueLIPCON0VEy8V
zdYkE1G/+qBp0USlZa7cJGnBr+B+tW/cUx374wHTA+aJ+jNtWIqRzT/UI9pvZo9n1VPTKSaAeAYO
ixXNlsnVRA+WdK5Ozbpj0SVB7+V5iiUiegq1c5KyJFax0/SS9RFSt93+5EHOk9GlvJKtorj4sElq
qTL+wFsDlANymgX+l7SBCIRwwrmuJy4/ENfVu4OL9eX3m4a9oacx4JRwzSyMpuyMDZsxHu+hntQ0
Rc3J9kFEdRGVpvFhYjf9lbkvpk2HkMIw4qtgrk0Np/Qo0Hf29skueP7w9eNjCgmVVXDTbfo9u8V5
mTpBEWhG3CnKJnochS6VRAa8N3XizsJT+GqnzFQ3HwisdCMMD5QN5yXp7yyipED56rQK1Z8nwnGw
Qgu3de85dq9Wl5TLV4RKUwLcctYIxZbt+VSjefSqKDnSBxQ5aF7CU2AoepLKXiTk5bfxkG5gx36U
/2reLR6phTsSqx0AoV4TAnWnTNh0mcnDCYEL77VUzsAEj3qMOCC59evYHLpgV/9V/QlNyo/yCcmL
vu53AZE5W57R2FPQXfyEzHQJcesGwP1lCtT36IT3/0l6ZKZG+MID2+p/Cnwk7Lbz3q3rRVaobp8P
FqH/G4bFDAIfAwPwMin1yoo6t8RUlR0N+dY7enpRgcSV6qbBEWlSCtDiK6wy46btbYLb+s3QpEz0
/Yra6lftObEGmoHsEewpv36EJmxt7nogRK34tEMuppnw+fS4x+0rorydVE40SUDxBcesZj1YO+l2
FFYwq9xAQHzUeDMbrD04Pdbk/duJGbi+8luSW3397G6JyWglhEU24Meq0mj7sURZgZIX+A7+7FeF
7q+ves9UTYHeYC8n1V0TYD66usf7cqzO1Hj6WRNjV+221wRVrLqd52Jt+7Lbl+lF1/SnSUss99TM
pH6mV3ivG+tEg3f+RhouOV6zzMHjUVomRVNER6754eV/DOSdCwgSiDfeE6GStgBl7mLwtqWXXk9w
Spmf4mQMcVY88gKPm1pPeXWB7pSzVp2U3Z4RNNb3pRWpOjiJmCPW3nboR/ijM+FTHfpZuOrMP2fu
XFpl+Des2/bQjkQj7zICgmQWj/gePJQsz4kVKyUwBQbdjmA1hlal3o8u4YB9kVbofiJqRR3z4fek
/dPujPoggWHvBNZYcWwnHC1plARYuqKBc1ZkzRkOBOzwsSyKZBl168OehZ1kpGU+jxc3gX5DNROF
vgxwav2HfAUfunsrZZJCsIS7Mynzzj7f+Y0Vp/3kjiNduT5CIH6pvrq5BNmu6pRbBZFq3XwTJPr1
aYeZ/RCx4elg9E+nWsCnWR5TodMVrpbTIese2YiQBsCV6u0PaJ6zO5O5wqWIRkw+aTMQLXsKKhSH
Xv1OWapI5iJ+O4kKFU14jed55o+w2iYIvYvcy8+/7JYAAGopwq8yJXKxA4VshjlvcEvX+pBG2ymc
6jL4gsJV1cjqgOGOmX1Yh49iZL/lv0HuzLcwXvAf0YkFPLDfFJljkEHG37xs4okPci/D/OsJ4uhI
wQn7upA06hwZz76s39tvJBS3+PuieLAZ1nxdbUb1yy9Uc1N3ISIiivHDtBBC+ptopzGaLVLrBAID
d5YhcN/PJKvnRdh1VZYNwHYAnrfh7pEZq262U6DnFLbq+vdjQBlQXU7R1ppieHZ6ICBPOrgIp9uC
lDUOu9QKTJLDe4aBcJ9mwhTOJmezaHmra2iawG56vDD2OVG+4xpAiGSfG9znVpRhQRHZYUTBJe7K
FBU0jq4UlLQkPUXLLQq9zgPQLi3pXwCjPV0TCoiyLt+u8+Gs+ajXWNZLvOvOBa4ihZh6qblkcFw8
7W7LcdG2OLzUzL/rNO45scwyCFKKRYrmJN3+CHyFgvsbDC3/eW5LOne1L6m429fozmpZPYyeLEtY
8HgIKDIK/t+iPcT8TkloFtZWDdkjN/WMjs4qvqF9/byJ+feAdInW0XuK0wdRxHSJ+1nKOGSRVz76
hsWNKDHx7Ogz7si73e5jy5lsxAYv//lvUvPAvOb13yodfT1jj3/JmdsjaIk8rPI7IpROJ5J2a+bO
fmEY8ccn4NYrALN1SUeYCfp8EKgzJbKdGCoypqSZaeHz9ZN5AqO7CNTdsdW5napFrCdiYxRslt+L
oAxnJVjfM9qvHBdy/xVLiC71kRJh+HAAqgttdAwBkTOmEpJP8NsIHqGnqhmPl5lXpYP8jPhLl5El
JW4pLa2PV+3h+J5fOXGuAyrKUAsZ7Y72aPjHOW6mcDcT+MU2Gmthp14puebijuaPvhMXylvG7aOt
WRzJ4Pq/gVSHMDP0KyVlsjKOqI+AwrNVDFm1vkZsVayb0uAZafRNHaCndFxCvOF7iv+igOujN3HB
mNe0K4ccGpJYY83lcosjN//9+yxl1+m8f5XwVIA6yOwR42eZ8YasCq/aPquxPOTE1VmLVTHJRKJe
CfNEExzg2gL6T3FjoDM+OhYXEagtAjt8ntNi5fRiLNGLwMLCHmYozFNAfxxM6oOp2KOwoYXerS+4
aqQIv9dopWS7h0eav4HjMtfcYNPWyofN2CH30UuC/9HEF9N1t2/8Vu1e0ZuxUp3OteQBCCNElbdO
/nCYiSg9U4lRdXJyjXsFwxpxBvn6vEBK8OozNYE5Cr+deqg4DobgCNnYtqlrEpWS1c3hqLxMsq8M
mgAo90rdYtJ38a39C0xyn2JbjOFv3lAGQcBVlvJ3T4ddObtAIaCbCcG5WbUVBvfTeJ+nWAqMGRck
+JW/UmOJWiYCki+qOUmcj2UoxYtN3LwWNtx2s3+YldXC5sptWNZ+F60EF0oQAAu1oa7IDlzc6kZh
2fcNjWmAer2FI5E2ZbyMSv3wBzqDzHjhrJJ42Rlo1l7ImAU1Y0smdGsnXxLtgnq2dJNOnhrezyxa
V8lhF57pNmVDNG8XxVCO4IDqaYdqwdqMoFVTKVm/lS2c+7OiotGyqZ5vQycwXsDtzEf4+y5cce8u
nx9H6vRbnAyYFG/tdud4QAtZ/wWVjSUrPhEbJiyMDWl+Q6Q3MxQCRal1lUAIMazGYWFYbGH0cOml
Aq6nwr04jzXYb9CeQumAMAp7YAoP5ifc7+OPQ6Ex6QqXYxr6VUCL4k4bOkiLYWGBnjiZQvztl4Ge
TwaxxX441DZechuQtc9g15m0XEfRqUem4KQdk2OTDQebFICQn62pz8Km+Drd/beL4wtb7eRMXzVb
DSzE3ocKlOW3GvSr4ccQ/ruEILv7BErK8wac1HdF7mfZgX5VPLl4eMHMcQNP02l8eGUY+rwgaUqy
rtSpytlj/hradqVjjnvswP2tQW6uFBVkwkxlDhPA9R4pQ4XSiWS3ecTc7pSYiOxBoD3RSjIE5Esy
AA2wofpOdBb5FUqCT+mXJvl/z4o3FvE5I6xKxalm8ZS9VLJXGo5nJ400lgvaoyiWvOkHAbtAJofP
LkCgJIZiBRK36zcPc9NKNp9Snzqy/mEOqUj5krfQLcIjuLw9byb/L9FNRxBj3PdE+IWwHqUjnvrM
YNwxsCyDnRtUEqFkJezW5til68+UKSloPRru2jpeMwbL9UXWE6zJkH/+ROdf4UtTeUVqmwnQPmEq
L9kmbinWU0BkSpRXiVXhHqz9C43tvOFAsP/By4PJTSmzvFo88fGmfaAqu5DbYbP8HAfLVTuh3rwf
Sj1CyWBXbfNGAASh2Z9slvSoL6gXohKQFVnFmWZ3AHW+T5acFLDfnjiFgJ57E6/NcYDitaCCb647
R5acnRrPtQqyEWhdZnLXK5K+Veji51IwH8zxHvEvlhw5MnS0cAFNGi3bCSdJ/o0I+dv95YkksBlT
si7AAp1cA/TSQElPMEpWtz/gAMVt+NPdRnp7DVqFejBjy32hu6etxNHFN3pSGmcO9zczLPpQIcn+
+6ohWp5g22ZOb0MxukSmx1U0lt0wMPkvZae+FRLNM+EmNeElMpRRQQLpDIFe00MgpBsGZAm3t0vC
5s4IRShEaSAtotOORJiKjRIL7uhZ4V32CorRUYTSbuVaa0lM7hm1yTcd6E8jdrnNWXVgAYypwcCE
TIO6hyGoV9QZj+d3s/KgcsrOVkPRWB3XfLtd3BkGfBdzThs3Xz2jLJ+/gQ+dASzrQlHjBQQ5P3Lw
3lZ+sRHzGTxJKZZB/73HwD3HCNjfSKlSmrIyEtWdmEAyQ5Wln+joPhdzXPIOhvPtBSQ79DFH6UmD
bp13kvXPcPf8CP+gtvy20hLh+tGiySzM9N1iar+GB1BCdrga2KjBzbCpuuFxTkBImsd44Nkdrzuw
RPB4/SC6ANKKFVWKdF7Wmrfofw8WPryCOMog7UClJb1KfyEymZAcNOhnfjkqdhL1D+TDtHk4Jdsb
2tsJ93qaI9Y08QH81z+q+q0QscRdCLfpIAAPek+GqKBqaOXIAgOZXG0dCniNB+7KvrF7rQe9J8Xe
ospONdAYgK9mtHHf80FCjwFwXi+LyWosr/nHiaB5SMQFvG7t+wWdLh3066tWqUM8UZjcX299aY9/
q20fwaGcbZva/yweAbvs6v9FZX4YWAXXpRsOifEkrQeg4kJ9p6K5ptM1W7fx+U7FZUVAc+cY8TO+
fVj2+BM/CtVv4iuWbNCNyLGcNoGSiwsLNfKnLNmtAICcCjGgcNBxqA8iis7E/WF6/b+5FUqb3RVW
9IVS68bYhgz1yU96VVghV3ukxQDzVSM2IcIoB+LpO6EqDdqO7QYFfaQ39r45eEeuONxSuE3zBRgU
be0J3lw3vNbq5Pfm7atLrKUAYnE35RjbC1m3eawFrT2r4zskCVjcrf4do28Tto0jo5pNjWRVYuas
24zxfu16vUQ8BaI87wrghiP/sNPsirFat3MnfzwuTv+GD7gX9nmmCgU2sVJHoN+s3dFd5Ivn9/6i
hBseht0A1PRWBUmXXT6OnukqjSvkRnd30edadg1x8jiIigRBWIWF13CH+x/tOC3fg/Mt2XjaBvMR
vJm063b/mzDPNC6JfwcIgJ/jM44DpRjZBxwccAwd+I9eDi5bEjiS/LXau65uV5ByWmXjVUSUCavS
6OPXqpON9CBRYNkfhvuLYLrIGB+zTWCtSn+kffNiK4g6Iah5NKyMNqOQEoAPjodXJruSIG7KWygI
sJW18/nYwvJ43VUE2C1VbqrPVKZcvErIGJVuux/od6y2Bei7HixQ/Y5DDZq7aFRJAHjLUtZe95NV
FH2iIafVFAWV9HcezZ/F0dH2l4/8TPMSmKdJ6vB5+b5MHH5krhgjm3ifkvQlm3oGv4k9i1a6whtm
+O77WyBZig+NchnYYfXA62T5zOevhwrsWAPGlx5m5nsgO1amFmuFxB5zdTAyGWr2qV7K8GZtJuv6
x/Br+y3MQV7ObHf1RaDAiuLtSnHbUrp8ZfAiVhBfwGmxWWKlJH5IJlF8XMo07jouLwRY5rANt1cZ
HEjfipC2mWpQdBdXobJwu3iXk0UesOTOXQEO4J8keV8BsFl8gFeTiTYGmPj9gkCz6Z8KbFDFeXz0
KOrSFOMBxhyVHHrwnnFeVcp4VhV8zJt8aRwWqaaKK2LaHA95Xv05xSnfBfsTdW/NRUc4jvWQPjT+
qn06OP5hAxuF5EIQeGogImRgrlP3aw/N0wpqDezMDzNGYZqOcHy3FhofYU9djeExm34LQ+crvoql
m+oCZtkvWnFx+jfm58URSueIVp9U+EAxqej5sa9+ZUOGQ8XNAE9yFRdYzpIK2v49U/qXfkvV+cW8
Z7kiIJMBLHS33KwaS0Q+JbE0x00d6o+Tg9k67Fn0dl59RBDgzOpYRUHSSHFPgKlZ+6NP77s42WFi
UCIevMQyErnIMCpqq9urp+0OTMsMqCgsljQoeveKfq5YrnfqSSVSaxolVbA9gVXFUBdsf9s114tV
sD4Paw1iBaw8qJ4z9VYAWwcHH3vG34uh+n7ngr18BIVuzCuqF3Jkexdc0TsdkkwsNxXEKguDCtG2
lKKKr6hcEnRKeuyVmfLQwWuOCW9VIxYhrp13wGTRSgEUsKyyTq+C0gz+ZR3V4vniFnKdE9zU1Vht
jJjK/m+nJH+bU4yKs3fxioEFyTXnVtr9aKMgVdTYNN0H6hmiLYKgA/De67TteMht2fpqaSet1HV7
e2O9NC0vwddUdVs5Y8t3eJi2qMm7EbG4ww4yhyX+AzE8muEwUe2ohH5p5YAK320CgZ4nnK6FROTj
03Dr2UGoHeO4e+FBafZ9pDPx8ncLOAIzRJfm9jD9if/hevJdXndvn4wlL70xSGx/CpVc2ZzeWM5E
XzGJKTydTfM/Z2Uv9hBzvQePMU3v4fycUIsLbpz6XXFBZ3pi+wuwJ+1JBsNKlJOID+PX06bPV+mN
drnzM/BXGW1ZPcIpbrRWw/Zu/8mylBBUmRHzwY5FrAMIk+33+NFejL9qYYveFovSg3uhUrL+9o6E
DQE/gj3t9iXiZnysn+YNy6p51S7KdYePnEKFG2vrVp9bC6ZcSAbTnKcu36DUkFvYpRaqFyisPGfQ
pQ48AsvvJ/I+caLGd7C+Eq2irfsvhENQvNdgwplMlPmTqPDoSsdYLXaBVG9WtUdevL0/5SAC/W4E
tasln8x1BQMtPVoi4X+74AvbjU/gcM/saq/nk3EQWsYHGlSZ6WP81XsMflQU+8J4vhIxr31BZzLK
8qCucAqES51QC3ngi5GfNHnNPtZkWC2NkjGdAPdKbsU+Pq+uW46/ykj2j9NnqxGRlKc8Pzq9Pa9m
Qrji6sglyoB4Wtf9y9HCQw77MlFnQ0wyUYguCoBwS4KNs5QhAL2OiUMYGV2y9Xjdz3dyEcrxNetE
Op3Oosf7QNZoupGFKsqqHBL00NjrtKiF0h3Xntt2OSD2ZQbgzf2fjySlIrc3NDQLtkqIWgcyMvM1
AOfwUPxqhqh0fboQGPii9wGZpV2rq8iUI/ZFBwhMSyvhO+XPKx9Ce/3nxLVFS4KLDaYGc0T9JPLS
Nn1o5YXzXan3RMy106812w0ZBSQZmHid4Oj4TnDm6xYlXJrM0CUOVKW/i9wNKBc5IEbzySwr778Z
qKmjOcBOX5rjIqxm6veH+53ppuNXZ70s18RXt/SMwxRIJ7BMZTxm0ZuddVZxf2BkgmZhYP8lHOj7
cvj9On2Azj8LTQbdyKJfXiSX8/Y4miJD7AoksHvQ/QkzliNQ6NHhXqbReHYvoeR7UhkyRm7FIDdS
y4x1TBTxLQI4lWbyLWH6K14KwUf3HZFOuBJv5vdeAUMohytPQzdqmCJKbhUpBbeMFvvpv/dk4A8x
unCdWkgwFOTLWCDuRrATvYiryEEwFE4XyYAqUaHpNlwyAkZUM8bV7JqBco6i/7jIzO7ACMlxrM+J
IulalE7tIlCXAKzKc5fEKAlXauomPw6w70A8GcN5XkhesJn7E5l79AtfHNqNRp65MSs1ZucwXVd+
18FE46EJxck1cwjWOqpIi+SrbGcTpzfhM5BRSSMiLdQ12uWvXIyVKSgd9CNLn73qJx3AVcW8TKW4
AW0MycPyG2CyodOTBrHp90gqZ0ZujACjXKOPA43zRVK8HJ1lbK826Tv0AIhY7otbmRmCfZTydyO7
8j8twwIh/33O+2gk7LiIBHiKMI7WAUAeMV04Hj74LmbnAPAqEkMB7WBRgDmX5rkLei/Bcoyd78H5
Kdj+4338akma3snYTj8oOQQPMJinyg3bDonT7cGVqmWGOsZy07cPPDADeOEl4YOO7wTcJAf/fKFG
mb2Y1tMH7/Fbv4Z+xTGwMtAd4JHhslKw4nNnO6b0/4f7Eq66/V4SDALhBaNMzk9NDNVUZiipdciJ
zki5WirJDIPv3ZryPr8DNjrdzlTa/9jPFju1QkVFaPgLmArhp5hIIqx6A8yg8L0LmKyMIQjeIPbu
B6ac6Nc9KQxCmIN9sBDa+cEWQkgrI0Ym0fGRiA2XwfF3IIuZWCb8AgbWjli2phily5FZUK0D0iwC
+Zat0rav+UjmCPqp0DyRjAAa1lNdd9kl/eghUrkTUSsFFPgKecNVWHFb9fgN9RkGYqOjmiwtfMR5
HUlhlGIWMh0HAcl7cpdipEt3D8Y8DfHrC5GYK5TsKhnNWKkPTU1CWq8IE4d+HJCQkHmLoIB3qMUi
TXo0CR6r/VMNe1t1od8nko/Dh9AEI2xY6+HOCG/RAx6kDTtg8OgjZe4AiDOVATv54tH0atRREobW
9XfYVzbizEJ4fqLTG4dSWU5uwiabjMrRBYxdSLySVzRUwHktjNFjVWYJg2U7TrDpXPFKZ/YKHlWu
dP0JZITgqBlXvrh/U34cbj2eZo9jrKbxVjoas0ZcLdwWuK2fEDdc4FTiRfxCpw2Ck/o5YUfDf8UK
ba/qChI2iLTqR3pG4wD23vA6QQ/kUi9HrXZ1liKY+vOXQWAjoYQ3oiBMWeBRaaYABlcs+MGMt27F
LovI6v3EE2jKsdKKMVOKRZ1o0PIoMsNFrntStvwCMloqGdTuZbA/178ROgqlUpPdqWfh9pEG7KgL
FUC0nD+A9WEpU6d12CLYF3VU5nmTVu2SBeorEztM97QbN9RnZCGz802Z3KcT0Ba6vvRU9SPCKNyC
BoU8vYnQI4VaXUgV5V+JJh5oCEfWTVYDnahAo+/y8V9yn9Xxf1Lk0mf2orE7kkPNGrxm1pAsy8kp
Z1fyKH5BQMF/TzDu/A95XeLKjJY6NHxJ073fUafo7RQdjbBkdNw0YW1MTNmVffBKC3OZDlbVmGgC
gyEHRWQGTWWPCJ+eOJtygbTQDp8Onc83gFQtAxnipwwbbmG2EN5pfJCVZNPKcFauZBce5mG5qL8e
Fh1tWtBC2QKACnl2GlFPh4zFhaZxU6W5TCzTVy8DreND3rnf2t29neDnSbVMXSIXGzd8mnCrN/lG
5Sa4vAKul27nbTQd2tTFCGVbQuhAAcdeOpYeCUWWelaGOUDJuVuY8/279LaCnwa3P55f6KkygPZP
0cZbpu7A/gVD2wpEtFMoSv20gn3GMYkfZAzOFc4W10Fy38bPy8WjJ5XEzFVsI39TV1D38bUrHIY8
9lywPWbxRsbTWZKwqVDTpM8U+/tl0pgu9K5FseHrgUI3LhFHkHVYBL1ZuDcZOGiwGo8bz/FDBOg8
aBvxrS5T/ukMEXhNNIpwSeKQOlyt7qXw9InFzBDvJgfKTrWYfyOsGMpc6x3YYru4XOv15kipFlW/
r/innykj7lBhW63LFTrDYtx8UbKgHYS/PeF185HEr46ZDW5hfhK62c3l4xyTO76y3jJULcyNnG5r
RT0qKlJHbRKyDJOmquhg9O+EbNk2p/8mteaJ66xQihsjU7upM1NgG7wmztm2WrmS5xrh6rYOCvxl
Q0XcJl8tNQAdkFMum+P3NqMhJPj2YwRnRN1btJiwluTW7JKX4ZoH091NtMbwgxlj2mQiIRNVkdH/
jAuy2soiio18AqJNkOpG+P6+KITp56LAh1GXDF8cQBQ9xEWpjw40gs3nr1rN0k8v9nnd1Dke1OJR
FPIEmAvXF6Y690R08ry2c6iGc5k1vpJifs8BKS2e+V0VShHF22w6X4XXns8mMYI/40i4y8H0+1Fn
S43D8m73SYFjSRZOLiKSMpE5n9W4NCylUh0oQDVvmYr9WbVdyTkqifVKlqp2g5B8Z2wSo+VtJeIR
59x+Ze8qqOpWVuXhZSheViQG3QjyypPMslgvpYJ9qKHYdu+WyUhuXDhD5UW/GV+BoVdOtDoPXivf
/kzMleXfqYIwHYwzdeXTVs8CYJcYooVUzD1nMdVzha5HEs3Ff6t6NKinFP7paM5zKJt9QCtURfXf
yHRP/Mg6ZSOiaNl+m5eirIKinoACEe/VKijsL2doxm5n9se1CpE/yxm6tNBgwy8vMvzFES4Pz0pr
iwJJUyQkVzfPFa3JlpgKw/RrW2YoudrS3Vs/fXfr09RMtcO142vAyJtZTsVsFNnpIivWz6rPyOhz
3sjcvHykNArWek74je4kcmmYosJPYYIjplAPeFQzvVrPZteFavdAEH0Dc193UAbVEBpBtb2lQCdL
jvaJvTkwlYTc52D/ULQq2LaWZCxGAgkj6lxZ7CHHZX5FfB4wo74/2cvGmQvcNx5FmectjJaaPAQ1
/nI04ljEYlTkNRyLPeqKUoi17QQyzlbyOI7WDza/a61QcSRWfU9edMK7rhijx+fDdIYPkhPZ9nIN
Iqe647vk24bhMuV70FLTaMqjmPkddOIb8GIlRx1iRHYGEPkgkHPZgN2ExfAGs5B/ozpkKk1s8V/i
ah8fd7CmA+FnqAssL/XSm6G2WTl/SsWX5zPSMjhkW0UpjSlm/e6d2pVSIDLsJEbYMXNG76uHoPJq
jreNordpFUls18R0KhBO3r5PDDmgyhYv6UldufNkjnAblbuX8GxlZk0ipkSINzzjks+yO76bIHz2
dXkupJ6exgtvC9P1iyieC8lPJl+dLlE+Me8biRUQ7/q9ybtJP1657LRHks+YiGPDpovO+CkspTdQ
7U8SyVjZ0sac2gDD0PlPGCWZWXkQwu2vJ3mYJPDRmlNYYxhQvWdkUCB23tyr9BLU6WXI5MsnmGLI
s+uZeNUhxxF8UZkWA4stqoP3f5aR3lq6vNRSqHEt5bmIid30EABsV18DeM1nkDbbCx+8+ClWruCi
B/l+G/k3yoaBuoUoHKPnT1apa5z8zRi55hhkDftbDSkeapkBk+JWyZ/HeyLckwvYoC6rK1QmzorF
CSRJ9njrYSgkLXxLqlBmrkvcPTjK9GrTicA9dVdcvDulxmWwhAc/ZQyysaXubDXZZC/imNRSVJ0K
GljcWjxgWBzRKxCRDMo2eod6DCtY2W53EsYmCwsyqMXGuyGbFfjTC2424DBCv4VAbgINbCkSIII2
PcQTdBcoyVSdfruViQhxZb94u/aa7rRvNPH5fQttP3P/R9jmBUf1AOVMFdP2e+il9s/qJ9FjHNs9
jGtpFKI8ftwcu3K0FY+SmX8QrqXmywU1KYysTDMa//1LhV4MXbUBEtZlaPRsRGBFd3YFLd6Dyvjb
vSQNuS7NRZuWfVeuU9t2u9Ri2ZgMCGFXplAP0cOUJT99fEAdwUzI54MwidZ7SPeAdHE+CDf8Bu9V
VmGaGI3iH7ZmEyu/OkxScNjgpkIDOsD20vemN20MS419Wmg/W7Ezdc+hyF11Bg+xpEZurFjukRiN
6fSN/yDmVtUTaTkeQA7hxYw01QN5Ql17xD5r85TSTkxnn0PS4MHN0cSqFBAapSdLMlR3a4qVoEvL
DxL2f+11MbXo74Ld1xIAfo3KNPVdm5P6doxSuBXlxYljC/BHNE3Vpgr2ohaL1AYFOWmlVJYAQBVY
xDg3AJTblmITIZs58nivhB3CgDGgfQG2YauL7kVJ7Y635/bX6uyvvZvyo8nQWuU0OE1fliz7XX4W
tJmjAjM40CxR/5CXMxTQA3dQWbuC9bubDe00fDc+ex/1fHoki8++Bj/oXjRatVjxRwwF1z9pHbLy
ec98Wyi9uNhSyNrvduTSY/zz88CyckwzrCKG0gWXoWaiAk5D/Dxe/Nc2soafcpkXTt/SRrvq1Gfs
gJNmKrVoe/66m2V/zf2Re7mnsXVePNKFCTHZ8AZa50zKLk8R3g1MjlOvAz0ykmtTxUOIBrXsychy
A2vhcXGDjCUlyHc2kTPx5JVjhqLXuQYI3ZqeAXNi2mK6TUCpB445lIkpV0ZlfW+W6jFrs0K1PobI
3nEVLwp/hWH7fOiRYK3RWWxvBXdfKLDxPdBI2KKNbEe87CIkNOPJOoQ5YllZ/+91MmOHjMbvx3e3
wkI6sI64PwirZSF/M0rox7Er9JFq+H3R/RKAhDOxHywWLFFxs/NmrjyVjZLO07sDhBYVrPWKFBB4
namrZFLGta2UzSeZVGMv98HgooAgb9F1SCWX/XJEm1sVjCrPN9ITiEPeMiRpWjrQSW4V3WDG9M22
Xd+azJAsmcuUBaKvLAkNoqJHFckIg1Zk28tcI+c7HwoTorYp7xc5s36kHbYMJQ/qXzMC2NxlZLWL
ObVIoq1Mh13Yrh7XigCsl4+uIjp61kt6aAwPpcwYCXInxPfUMoU5zpLvyW7xgpJ3vWQrNklrnSND
cigYxYtiT/ryJ/MmyOta/mCI8aNr5pWNpOqLbn4FYmKhzXCAvdGlj4r5YER3FBiZN2FIHGSJdbq2
c7pEm6l4NAiYsHx8O/a2fObtN/RDXbsO3dkC4dBnRN8+LhZE55CtC2ajSb+8svet0b0mrJp4/0xj
K7aZ28FUkKqoKBTY6RC0KK6gZsxI4Ex0iSwt1Pnxy5hAwY1UPw2/SEJs10Oe4BPsdSk8o1uKbK1C
ja8+ePRq9fNIG3Aw3UiYcklzDWIkzroQTaKk0C9JUSnjiqTgSK7LRST5DpJhtMSkr4mCkWuMaaDd
vSHIGXwCBOPgqKuunnhwFoNgctJ8+5lo5Y0sT+GR3YnorEantkDFuXprAzeKSF4+tbjXzLnwQMoN
zL4gTq78DRhb9ta6zorvbvQwhFAUEiwhGZmVQE1zQofuC1TSuSt3wesvuXKTpdkc6c6bojduH4Fl
XxL+98HaxcpxfTtnAhlCClm6JZi/OeMYMfBbpI/vA+odrCL9bxMeIOqo4muiThWsba9rvfA6B2Ll
9nMwi4FfHZu3y+D5C7fNG/f0KE4aHwGyTIGGixVshR0ls/8kQOU6ptLL5rBF9dNX3LXubOTlQYFZ
oZWIGecs+iMjqiCaAXKAT3rBliFLDrFURlCDPEd6rvTNfAhiPU8Iu24x8gJD0/pKFz/FvIv8hylt
bOl8jt9QRRVPiPQYg6ymUL8IGd2Kzz3fGVkbym5DkpGhm/7oUVnRhOCrE46BvKAdY1ZFXVvjLl2q
lx9EcNdyk6HvoUYqFyUN5KspZ1u90M6S19yTMJdWkfU2/y5X1t4rfRXCaQQVGnkqDe/6SxRNZ6Tk
Tuc7B3LT+DNjiGp0AoNkglYN3REpiCsHpN9FnEC6FXAuZ60gJUYO8KVPJ75JMtE7SSh6yTp5o+Ul
n/P5Dc0gOC1zg61hTWERHlHl4/Haa+msCCSuOub6/9BX5pfrMfuaGmTekzPhARIgEIOuYPnXpK/c
Jy2v5uf3XGlnjX2FcwzhnOGDEMEQpmAuOnc/mOmW5oJS0ZZ2kCnB/w+qsZSniVx2n9vHY8fX0M4m
DQWADgC0bWUj2sr4Fz8Ko3uSeTCx6j/2UpxiUOlnb+hnEkahwlwBfhKEHe9n2HwDaq/F4amR3UBL
9j+rIVIactfBEHS01AlNFPOmBclP0aIdWRiNVxhUX9YwMgTJUs7JlhMgQ93MxtvCOi+DQLUcmAs4
so8bCWWrSAZMPZF9v4U002WGbDBRHUOS9HiLhLNMdHSJQc9N+HvtUJX1YEJTbOALZLeVZD69z60/
iLsb5Ng7VuI+fO7QoDmKYg2LNlUyPBNTO8naXXe+Y/0pJPaI/JMYVKmys8rUDT5CU+yeeEWq0wzf
p0Wpm23yzmunYeH5WHJ8oZsZ6RzeIiJaFQTeuKlWwrO9tuM79nwUud2FNPvZivfEkuGJLqsUbrKD
rDDMNR+0+sJI7Z7c4AAM0XAIHDAvqV5Lln9DwO2hxbLhir45LOkf2n8cYeaJFVLNiX6BtsPdveV8
6I/TSRllRSTi78XaV48UhHVUuAt+/vpB8XE+vG+RhGRBncMI7XfX7G2kciv1MWmbbyh783yCkfCI
ECqkO13HY1F3rABO6ys5NKP3HHAk0F58Tvsb5W/p/ze1NcoEpa1j9Vm4/V/gfKCiOtwb1f262Bmm
6PayREwaByFAp9O8exOiwIbldQHCJ4F6qWsWTqayDjrIYbWCF1lNRYfnV5/qozpRyoITkEsepVwm
LV+TtrUZAlPql9BHyYjmTAar7HcR2Gao8hL3CFJvABU3A5QltQh5CpFg+12C+5R/m86uJsoL7wST
HvB4Ia1SIAD2uDstaBsxULjrtqRC/N+T026J9csRD7Il1L4dM3anRHQIGW0lt72Z/Sqtc6Tosp2e
2e7JXtb1+dt+KantzpVC3YwXSBUXwYbLA/aWF/VQMq464eEM+a+LrmVaoKrvN7OxYqAvFPpWmLmP
WzyCOvCdRAip4FVItoYq3f4Z2bIUmvRS6Vi81RXAFZPvWVCMLYioXLeUY76xnafRQp/aGg1GObLT
2XBPNAdwzl2//cPZ1HzutaacxLZJS8+KIZtNrNIAEn5kfGwwyR5Gyohr/APe9emg+jBWoitLZbIW
k2gskFcKscxdOAyJ+8TjxBeBTvrx8eUVhVVloLgSYZMbxTRaMOzJkca84VMU086pY2hLOu/3nxyp
C8fPbu02nmu5SjNs4TNoghlNukhJBPlcbQZElGVKKJ3KivRRCVIUlG45DEnKlm+4OG5XFbmlf7zx
id9csD0N73zYGwrmVLvFNbbSoc3A5Yb3oWzuvQj7vJZVTitBTA7QWWhYj6CUsMt7JqkzgqPwM21t
Ou03+TovqI+NnJL+cdFoR/0ZskfS+fdUyXwJoHFEYLlI4PGHya82ixJW0QaTE6VyELiDBGML0kzF
kCkvqGkRBHAuLDALp1R5+6IutEgIVOY7WIr1Fp+eGrp+9Ydzg+cH4xIy7ZzbQYyOqIck/I5xsQAz
o2cvX1UcPl1wGCdRg48eUC+Hl4hCTCS8JonmZrT39mb/7Lxu3V1W62fD/rEUBNcIyh+K7jYZBBJp
ky9Duw7CBBoThvgV20H3HKZkTpmVW3xgWiAEg+J+FzIEJciwn2rmkuxiEVP+F4cUOuNkp+Txbx9k
OWEq6oxKZAl+MeHuwiOHjqsm5uuOqrD/EDg6gXdWGPDZ+Bvi7Ef3/k3O1kvfIrqlUAeWuTandjiR
okLIjbAmAJRdgtkN2zX6SK+Bs9e+ZZlNPQJZPTpqdohmUORKjgG2lrXu3vTwFU/QSOwydK/p1mCV
0J4/V96VfTL6JZNZIOsyc1EQbwMHQxDKTIFmbNRPLgnrwHcI7OYE0jn3HysyXs8pQoKPNn48HclH
CVrcX9EsHhdYtZU1+Zf4ukj+Bj4X+l1uynOZdzpWjhv0im1Y9KaouPgP028tWllUU47mJ5KRCZOC
f1wvNZCy1u81YmnN/pyofap3yyPOlkbfq8P/mMEXgHzyPEXEc/9Q1QCq/HYuy4/Wsr82Rd3y03ZP
ZTHkb+BLmti4nkRTWu3m8BU+LzFN5BvFQhywxDrsRIVkd1alEWM+FoS5vU42UAgAoG4cm6n3LNU4
poiXQet+7reClwNTxHw8LYYwLvJUNuvJzkV9mC/OV7SbGpBH6WrVt8lnuy+KYdyeTX6Jyhxyau/c
rWEnZ8XTQIZQbczmedlzw8ClDcBjyjb1sq3ZWZ4vwy3EPvhLAyK436i3IbmBIeoiYdyPdqf2eanx
mBOW76lHSkgPdebEdtqVMuIy4tJHxIN7d9xTqE45DRcvD/LwQHXaFajxZP3LkdOuS0bKuViyVi/3
EiaCXwDrfo9LgMFlBj0xiaS3SLaJj8u7YG80+GULjH1/LZ0LKPH+qW+vAwYVyvv67oLuBnvE88w9
UmkQoakdSTcoO81jnvcash/bGLoQzEq7l8ogQYvUNr8gZv2gphVwqLKuZVmiDnjfBUUGxmjCK2vf
BYwCkbMX5FQtLycdmEMBUIQcJxqKKnUvwtqrKW7enjAXMUHUj5PHq3zClKHeY6OK0OW4a8adJ9HV
viM3puRrU4tmylS5Q3FguzFFIxXBR5PCYQGKe6jqwfbEoRtoE4/FPqwMGeh0D9HzdfDyeoLOJwA1
epMTFsm+lLNE0CfuMOusQci0WuFf3IPXYtR9PV8oGIybsy5X6g1fuMdAu9cKJ0/KbwZTSYb/XycP
dnR8mTle9E2VTLXLRxCSOpkK2OiEPDSQlE9ZcHY8YzvdXkro14aOlo0XwKYCnndn2J0OZluFUjwH
Kjxu+xwfr9EjLGmjSXsYQYftfJPj+14sqC4e0e+aKre1dbQQB4UFXSgRjg0csm6w2FmoCR2GdU4P
HhVv3gf7/ESdVq1N1gxEy9ZVBzpn9nOvqeu21lEJ9/w8g1mLcxi2S7knKhHuiT6TU7Yfq9ehihOF
tj+Bu/5JidMCrYdh+S7KfK/UkCYCVRyDqPx1jjeEF3dpp7Opl/b8Pknz7O++XYjepu2/t7Lggh3u
NQjFiIecL2uv92vLubVeJnmQoecoQU6xieU8KMc/i8pJG+ETgT65mb/TTdxgychvUXkJ1dzTcdMK
kes47sWw0l/8MlfsRaXILg30Pg06IiXHuTOCrjCBbGaSWIlZ1cGpGRnvcyHPylP4P7Qzg/H+ZRDJ
Bf79t7bGin7T1YSwBHhtsvXia8kaT0QwhBDGnJH+CiB/9jwdcTLvrXEqamyudw2wN7cZ7XZcqSk/
F7veGVwpiLD51tHbrpVpMrLAcG9irv9TAtpzb9Wm+EU2S3r0reSY1LS9xs8bsbmV7tZfMe3XBvC1
Osfox3ftLeSqvLlW5/Ku7AbKB6whVWLUN7h4knvG7XQooo/me+fe2BhPs594qXa4h0SJXCinT5R0
4gpm7g0vxLH9DdNYDsTnayq2Eyu2CTR3OOGR+uYkUU9YxCPHuGLA8WnEPB4x6Vte93X4RckX4Ntr
RlVbOn9Ryx74q5ejAxkNfR925kncJeAshMeBVAC8/yh2OqC7MCM0HFbQhY3BFxV4JB6CMtcFeu3w
twcjyTBKgE44EP5atcokx2dJbDNEg3ZgRVVdE2fX2Fkb9RFbJeV/cwrz2gwSM6xidoXTUKYw69KS
xt5cNLJqq9QK1/1F/0Fh/9nEv3D5LCyTuZwp7C5zX5UKww7wzKfHNWumafI1WsLUjdbt7d/EfSr+
euvpiSLw9sj7q1Jz3Hc6Y29L7/XGv7/VuuMaLqU1jdn/BJ9CzfdEmVeDOapfiWB5++QCMHqGkZXh
YB7EluAr/rsgzRqnZQaQkG8EVA0lCQP2cJ6TNhQa+sjXdYbBq+zVkAVGGN1wdlxO9CkmZpceEoyZ
1B5+OB86tXVTW2cq1xXDgV0Q6WMqcZQW2GkkL3LmG27gvdW7hsrQ4zmgr7zCTa4X1Ui3G5zxI0lc
3esQS7sZmzkfHdKQ+RuwdDbno0Mrs3ViINCVFIaNKWBtiWucEIctYdqySMOXqSYNcbsEoJqC26iO
6bBSuFR5DrR7YUZf0cB3Sbr5zLXk1sTJH31IR87fxxt4s19zThL0kOpXPXEpVG4obskwz0jy6yFI
/Ee4kTOPeGAW2smTkP1O0BK7lQ4fFN67LisDFzRntX56p8q9qaZTUa/okln9H8A9vb+InPvYoTsb
PGYNGYewnuw2r8GhMFXFa158ZfiyHCelglLjWool692YCMBFWtnUiujcHuJzPqyjbFObFFiTf2dv
vdr57sqA+cA3opwyTRrqHPgDIsbB7cTz7qJcbVQ+UQgrk9QlVf1Lk6Ay/BPtniOMK+XZVOPxOh3e
jUdk11ny7UtfPk1szcWgQaCPDe9oKooBIKy5pVYVcYU/yzEQiVUZT2hYe2tkg0GNYqha/TvhRcPc
PZrFOi+h5qkxmXa4lSsLcP2E4tQoMvLFsL9itVOxyiqkiTByTVCG4VlHG0J3fYkcsexr1GfMlpyp
E0Zh1/K3jNq3hRj8QagxpLdYTqtvq0HouJPJP/tPfluNOs2+3E0JstavbT1octQL4H9Cof5NGmeQ
DLBNrAIM/vtq304qdNzD1GOvU1Q8NyuqgZ/b4soPScaCKA96EUsTy8U2ROBlq7Rd2VRM3g7twg4z
oF2e69kmviXzWIpee8dHCsNdR40vIt1qi+VuzRgQJizCOnhj+T5ljWBc7YqfbFLBwJfHyvVVgKqX
86urjvoocnZ8DRDwv+OwTQT0rUoXwVfbIaV0LKazd8UfaDF+oaUtiMRx1xfAA2eQ+U0eSaLO2LGG
cQXzhnqBKbzISSRuC9T5XD+H/aiLM1L0qfHo5af/0/Hab46aF18o5XJE0ZN0ES0QryhxLkxG+LOL
TsLxyHhCkaMCVP8rNxLo/IKjDlwx6dEbD2+QbchCKCieX+yJiOMWXUysPSaWTSwC+X7omY5Z3i3G
KJ585OpI4AW395Oh1FJWSMWqTnPDWKMBnFRm26ieBvJ3upqh0lF7NM4pse9ESacMhbmEzNdhykRA
J2LPP3cywgBC3k7W6nd1mDkuMK0f/sa2FIYUc4GWkkhDmQWx1BAl5zF/b5BFbh9NyH8J7V8iOLn8
MC1RGmaoLZPyWzblwfuxdNdFDMZQR3WEnfFMbaZC/SlF4iC1WOoRwotpoHs4kuRjgf3Xiykrbqlo
jTab6iUpeNb92oagDc+aNZytXQZ8/2R7gTIFju8hNVywxiyrXjjC4lNEiCfmut+3ou7g76U4L3zv
Q9QOvyHiQj7Ldh6A0Vj3llLbx2QqKW7xXb13ejV4itUptt3UMZtSBGpV1x6ulAUtf4p7b6o/mhcx
Vu4HrASJH38URbDRp4PFPFXtlwjrgkgu792534SHnlinbyIJ3WywsaL2ivS5Qht5miG9xyCulN2l
N3wdPoDWhpzI0RBRAmYUBt6Bej5EIdwfabPnqsJEtQLI0xgMua4Xy6cwkKX8vaFFEdjNTZCIhPxO
f3HJiCLKz/fmk2uxQmda6ksXBDpw6m4iKEwr+PyVFL7uFHdJcbrGLdoyrJHGipCwP9ySqnHQiSPq
PlKMbnfEDo44uKdBDiuODT4j8cEkxIJpQ3FgJnxHSGD8AE+tPfSe8GWWl1miBGmKISRL1ilB+HFB
Pp7VLXMBGqI46hV3jr5IZiTp34D83U0tEF3jbG99ls62wcEnfTNRAnVtMyAXh7fR+u/62FXHEmhW
2+m7y5N9+oPWBnGpQyJaKAzl8EVScztb1EGHWl3vi3tIkrTDwzdFlMew220XUwxlWCsBEBEoXGtd
v2PB30TbtD0+QiwB0YZoj6CoUGPB1JB6RzCPVDyHB8nI/m10kyd6RK3574zN/PTGnVDHV0o8kcsd
vqwrd40mhYG0WywBBhQfg+rD+7uQPzBBO1oCF8qD4kKKTTEWArEgas82S0l7VXNcaKpX9bOnIdyZ
2Ych+BvU632YuEMBWxiQAX+jSopBGJvFVyazN5mx0L+QOkRZ4Xp8X72ffwPkoHN1bCT4x0Gzz6UO
hLRgR2ZeI6PxNISpCH/tJzpBWZGKtBts/cSZ7WqeO0lVVm1dosVBnZgMNISXMzsl3Q2p3H/pngo9
7nk3ymR/QEb4M6367J44d6hXzVDERxO4qXzuIGUrMJojcMfP1idZ7DbBQJG6VZdbUWIcH5yGpyiM
OKP+WY/0Xn12BK5KIQVI7BlBFmoNYfh+BbW/2zmphvvNuZUfNZVMnmFxjCu/jKGZanVq08URD0Qg
MT9O1jKS3Lf2DrNw7dhEQAIX7dHq5zlejw5zuwyoUzGDyrjAB4Hwl9Mh8kBqa0JvZvDi0ammYjWv
Nug4J69i5C6CkNoydVqqfHIs/rAMvdBgZNxQdV/n9viweIfEkKxxTB/QEyz21RVrx5luvzP/Nxu1
ddLFwuqpUoSNdrN3Tbswt12oEgDM9FtTplLr+fHRt4q1VTauFrPaR91HKfrFFhROExr1kB0CtBJJ
b6Gh4zDg5+nLLA99Fz2MDFw/vA1nZOFtyWhQBcSVpGT/gassnKPNyPY4mA4AB2/QtQj9COUW+94k
hMx18TZ8B6RhDgVXoyCpLo0quNgIx7ksOONMGsjrolIKL3yhH0lb/A0B1JkPXoC8A8TGrzuMqUBL
58A95trjKHQAW5jsdtqW+DbeNGbXA9cj4G0cELU+beSTwb6MKviEGOe9JX+oUvDvxZMAp9dk1RW0
ib82XLMiSHzxbiNBneYKp4/YIpSws9joVO/p965J1kpoi2NIZf9ISRbBygYyqtFRpeiH7SAOMO4g
18q5nBbdmuUzo9l0NWlM9yFqp5ysCAHLxHij1Kl5En4pplHyoMXCSCS1RNi7liIxsiRFpkQCHUkY
LM6nR3z00MBdQJQHx+5hPeASx9DBoZa7AMR6DY6h4ZfYfdUC/7cNmBpwUsAZPBPE0hRJIcpGwF+/
tUxjK4ep2ofryV//idH+UWKzyV2NOCCqkCZv5/HhYgt/osTFHuKXJhMJKfGWfSNfuEoJaSInw94W
AqA7mxZ6Lljm/M16brAA9Dbxgm6UnZfrAUTMIzsXeg6IGFjCC0GMSWcy6L5xNd9DYs/oDk5Gsrsm
u+1dbWQjmyklzMcNdGSq+34ggEXTC7gQcIMLx207HuXnFHCF+GAi0G//Nvamj+Q0HZ5Nj7P/KQ7u
ZRQMnTT7zad7+6cxLaUbgQhr1cvYG+meVvOxeum22pVisQjz5qehSws1nff+18DeeXJeJ42XIFx0
3+s83kUoy9O2nPijQln/Jj+5JQsDAmhX/6vlKHmV0l9IV6qTBan3LSBWp9mj7t6Ik6Pyen7gUC6a
M7NA1fsRWlYTk5tF62qduJf1MX/YWRtyoARs5uha5KXcvWQoqS3wcGS7P6p+nKpawosv9EdcT74S
UUsryl+3RVY3rk3eqUO86E4LMMmxprMIQAmwwP5/F5ShDEIecAxYkfAOhFxDu0SN5bjYeI8me6S8
O3DjrYKgeJ9YuQk0UmJeeK3P4meLJZinlSYv5aEjWCBRAfBC06qcQv1LNbGbqa/gVVoZybIHSrR4
fUV422HaOb7JUlVHRClilsj8Vb01au9N+G2uN4zPdxkbihst6MlnvmTijUiSTo3XAs12JnapAgDQ
SqwHYMbOTJMvQp/ROAzlqKHzKX54TpRo5XDYn3dK3Wn7wgPwpc29k2DRWl88TcQnEuf0LRdKQxPd
BpioqldRnbRIa7S3kz4+AMUG78UDuTwtYdbWQAMQzj0vxeLQREVrLnP/TQpsJ3V8/ZaY3GLqtoaV
0SEKYAorMSeDQITqNjUZ++tFtE8Pw+KmNj7GVWbt10Vc6GMGrG4KjxPtwSQeNaoBFqX2WcLgCk90
iGSCKp8VBR6EwVPTdBjeboIfwzWN4vxWAFXE5del/WPd9wCr9OJd+KHdv/cMo2EJbdggt7F6sx6+
1DjvVKIVVYRcgcgk79Hpg50o1UT4DR/SPBjyap/BIXz3zXkpMwphMAhFSlyGJ+kgyHQGRC3t6Lqf
jErT9UJ88qtA/FKT8yFND4sek0vfi/iaqd9nk8qrT2feDshGCI7XKjw+X/Ph5JPBOutLSXCy4tud
sJF5Sc/nzdnxtqvFGlqbfpDhi8HkxwPQgOK2FWdGtTK+tXT4NT55FYVTEkmUoMNqSsxUa37rQXpv
ygqgEmatDCRvjt8ST0IMOB/6ENmv3q/rkjXso7qa6QTbEpsHZ3ui/WkP6+m0sJpQ+4qZbj4Z2hcc
3UjHrLpy4siW1dtKYmu17makI0U5T5thxihcVBQ/SiMXpFxgjZWSYqxcTpcQcjIQ8Ih5frxdzDvM
FMc33UMQXXV5DC2nqtYPLGEbPuYQtkASn17d6ygvNkbfDkAZHNGLAozEMPAmkNVMgnHGaUZS2rQI
FUEW3fghkexetqJrsPP33oX972ezfTZdRmm3NrUgpClYSX1ZEh3jT9f6DlS8aQR1LTUSIcWe7zAy
aopu4aEu1Z5OSNbKBGztekzgkFfTsyrmyvGc6z4PQ1WRx1Eb7f+P9n9PwY5/sgvOWe2abuzUNR1p
48rxxKiHZndyEMzr1wxnApdHQjeMc0fyy6eoi1Gu0OvdcwU3bm71OFw3TeMgtuqZIw8zGbTru8dY
l/B64dCcabBDDuNmoXnCdwlW2z3GdcEEVNoQpx4s6vj7BMxB6AnesAsMsPRBgDXgQs4IQHa2/JJA
8odbcueFFiZVjtPoT0+EDNBnUfE2JJnw+kspvwV44/WKxEod0Io6saxqFy0JxLTXIM2kKYX71ez7
mdDeAJH8aW91Oyu3ej8mLcnxnoW/PH5mQmmED6c26BCENG9hMIqITAM6K9UwPp1CVepocRe6Ny/8
qhr7AaVAo8EPPf2ovGFu5ViGrmmN7QZ3eW0OJ2R4gocoC8gzPgTrhqPq6vdu5lqgZPEn831AAspL
Erfw9jGLCjGKr9cRHJuDSkkIDn5qYIsYwS0TRmfV3/3dMkxcxE8z9L9LjtnJKsE46bXmciPoaYK3
O5FdYHBa1pzM+p8sVpqaSLwaTJ1UrEMeUNJLrzBDbNf0nndREt2BweTcxyR8Fy44Hq8wjV13it9E
QoaJOvt/YUiOkUbWPMJ4olAGPkDreXVlbkO6oUbFPc8+cH9clMUxVwVKLZrkz+7ddj9ob8PfFNi/
6B9/RKf5/vtZBadr8gOHkTjWUdmbIx/jrrQaVpx8rVBPVx4cZYVCwagXwF5DBgdtH55w12y/KUzo
5eCaA69nciRzvQifjGZpVmQoBqfKW8mY/7A0QaOUhXpXRc/Qsoyp0zFTS42UssSESn9CP5FxMhBW
831PQk/gpizOEcmVwKZMR6N3teZGb7CvWXtflggj7chUy5qyOWM/Ut0yiB5fAkMLUr7IoFATpk3p
ZGH0f/gkZ/4wSPE6PcgFPrkTWQ7x6iYXrBQU3IWwJC7kScQVZX1ySBEFBhiYfNIMs/sppxPV9iKy
LVANRYmtbY0Sv7lLoQaI1ACIlgKEJNx7YxVNaoKa7tx+1ZwIDM4yixpe+s7uW92E9WP9hxjSCSar
oQB8rBTzre2YPa++1iT/n92jQemy3gKHxS/1tGayA5FGmPw/9YX+SqUY9kccAqAMRBwDs+wVxmzr
Q7elHVxO/ysXJWn1LXSAL+YYVF89GW3VUSqExREoCQ/W9edPDmxUsP7dgSbOdacY6mRDrsaADxxz
wUhNw/5HwZrM5h7tkYPlastqM20UdNzmajWmeUkf4aL/0o9E6+NEdQRQwM3aLJhjPfldjuR1C+cN
aOIX/f8pj590e9gY2cjbjmOunsyGuy7JH3BUvwE7IR53/6y5JqcXRJk4tezpWUeloXOi4wXopScY
OWmaRKu3nKldWyQqTf8gvbnT/Y6DuxC/RtF8t7/kFh6de5MUfzab98neIvtvQ0OBo428Ky/QEIy2
sTe1TLYx5yCn9ctLD9JMAGA1NBMYjHDt2hp4zfabl9MfYPkCW9Tc/p2a7FkE8bzwq63FBrZqF2nr
9Isqk0EYp5hyTkARL7ApajenJVQ5iqqCOFlS+ipN31gmSabAiG7UG2GpNdaqy6JqK6t/+wFyq6bp
wBmV8ZvU+KwAyShSBUkFIt+J8OK2ijI5KcQvUkGutWF15Wbz2z0QFgEnetkx2wt8nwGhXFVNyWNt
UqDPexCGydruW/nZLba0TuWGl7StfdbNWjQwSjo/t4u6GC8fcwq3sCEa58j6bGkP6iSFZW3qlJjK
ObrHwsLW6SWV0QJNGO8jd+OLiEIvKKiL38g/qeVu4L47W69WDaDCWQy6NlU4X2nb0rl19uYb0QIg
PmTqV5N1wlJ4NtjwG7jR2O/V0XEzZU7f2Kl+Z4D1JPrYpQ+F6hwUDMs0glg7IHNNyx6kIS38dNaj
VNSftLfmivOdmHi4NBSkvHX0gBdqNiActAy38/viQFwX8idN7CMLNR2aJB7RciiiFD4pVzGYiQqV
fpIY+ypTgrIFmrWrx+hquZygIxAqueJZu0Z+BKwyKhItbDiNvIztPfB56YNlFOsCUddSWYIBObTH
gBbfkDLBOS5zjeIYLGp8Lp/+ZocRwt5WRhpbV80Ty6GtQUIsVtnckbf5p+iUQ+nGtYnOSAf/9AYz
hYY7epKcox2fcfjS9XImdRM2OrUylhZh5k17y65nceHfc2y8pGWvi7F0lVnvrWnUg2idrd/3LE6+
MVLXIxykWBMtf2tNAzqUFKXIP/gUN9JclFp0olgoNv/F0NPXitXJ/+D5o+HwNvoGBgNzA3Or2qct
E1VsyJoAVsaxOCs9R4DpsQR0/JFlIT6EFVDaG0ZkS0sbkqhCaFIr3yVqYzdBXCq1NILjMacEObEu
oZNBlTdWhQDJOlqUPNjwtr1NjivOqVg+kr3E06P0//yduTsudAKPYuhUL9HghsXGbLksbdJ7e2wE
2BnSTy8aZXvAjemdh4NROZEhcbuWufH0vsUBeHpO8lIpfBmu+ydhLSL4TxepJ2mTcTEkG0Qd1h8D
QxsysR9AXmFUECiJtEgOAeSJpopONtVtCNGVK4P66D/aWddjh1fg8J2W0Px1HUMEUV5hnGMUzjvD
Low+fHX9jmq/0JxSNp2bChkaPcO6/M8X0RIbnmeyc0YyuMiwRylo6M7VloU0jPgiGFcCAo2eskGg
zfE8NU1lXaZECi0w+iaDgf4b61b9BzXLlxwn+Ho8EBIzGHnjUAoNPOwHBKLikeCqtV0KZylnKwv7
taAZgxODnoD4nJbAwLI8mmF8Gybsx6TvJANCkkktGGBDmzx93w7Av/mV9WePm0Hj8UWNuXsZA3hm
T+SOyZTsv7yvFiXReHbSW2P0vJrOfwTqEOGmw6zkU5upCDHo6SWdv5GkwQiBUB9rvqLp5djDo19N
aKqUtyu2OLSCdowF3cnopYoPRYrn0fG3ELg5Fcj6BJtLryr3m8+fxJb0OcAKPeAOqW4gZ5pERvs0
xHmMAXNX6iW90Y+f9yvask5LQ9znotPsFN/v9mkHx+PvhwPKsGmoyIkd1Y+tXRjRrt7+a1ExpsF7
R3XyqdbZCCnO+GzlajM3pHoGCAAAlrG57By/KAnq6dJ9z3sa5w4T4m/+Jo65Cq5GXJ/LebG6/Kms
sJuE5l4WpJZ8bn3pQUP20zZQmci78ajPSKGMmtM/zFq6cz9rOgdpc6cTmg8mBEPwRYW86hKD6wGt
35qxiZzi8zV6Nbnol0O/4kBxFiBTCvYwT925iMKGIib08g5pf+c3nPTsAu6LZ7HbYhV1ZCblWyd5
AwaNZe0blkaaLNroA5y+9T7UL7jMkA2h5OGDR+rUXNOpLb6UDxMR8YdtiykSF+u3zjOKJ23mseoT
0sVp3tJ4yEMTRdzluNN0c8CB6JV4rgL+0yxR01cbVwS4GH+A32SgjpGrCP9Fo+737wl6dz2E4dEj
xyBlnBT+xImkh3sVCmDd2b4n6A0H4F/7P6PDki/TiGVEMoQdZGACR4rwT9w0tZFOvNpQpJGv2ufK
6kyiuU83+xQZJwhybw6BnX/heeWCPEJ8bHl/b8NRWRCNg1vDtScUd+/UD5XTCqFhcBo6QCEMYvJF
hHb7S7sHcTBpiroOCpopFAQt+ScKa+zBTHe0J5bEtYt4crs3bpWz8Nhr94JFkl9d6k1kffqpnb+h
DFIRMHJJsOi/bRsm88OhFpTE+kZmBlSXBfx1PsoWg+m1SZRYKh09mK30Vc5ozwKOI9sCxMaudVIX
u7+u0HlDCpkbJsL5heRG4nMtXiz2Jp49ys3dU/83vDrDouCZ14dtJ05OB2bsUQ3mC+i2Y1LhkAUg
MtU710mQAHd0XXjYtnuGNsmV/QkhYTzFcuqitvsPRjZVdk6JnS2nfoA3Mbtof6Zprv7dtxERIUM0
ljujThjnxt2qpji7GQZB1Di7jzJ13znV8R30WWUeuTnLniwbAGTCQ/dKFP6e5UrhSBlraurnXoxU
95rRYltmajiki/3N1WqiUmKSPqWmWC74ZHRfht1SUrbNYg9Wjw+XwrtkhTXglrveFKAATPExb1Zo
zvgUeOQa5tRWALkjgnNH3enFptkNub52kATlToJQWiQ5q8vY9fxOI85CBCk0eRq6hpYzxk/j+3+P
tlLpx4N4SgmxSew8Sfqpc+EVc/S6GadFRcnjls+wabgkU4ZllUDJKzABdyQzIKCVpbQgQ4y/qal8
OP2rtrKTVwexlSkS9XGYNmXWCmndGKFAOnbCwAcrjChDjfpH0hgYd2YNVL+AQHoQxYzWKcKdYQuz
3WhuqRoWCZoe62AujXxQieRfVbYdGp6SEetIVO6jcF+8mciPMz9DtCaSbGfeaZ8J7tmBZDaMnd0G
8n0iC6K0FDZ8mUaZxtrX8lfH9YlaebFfIQ/0lC3nr2BjoNpBVaYkux9TQBoJyx10uQkld3oeK+jv
rbdZpdxxImJsa8DZkowwM4QU5lyVA5TpKA5le8jxkvSo8SY+y8iNAaJ2Wuplbq3Gh6/CBq/5hre6
2mJWGVcNcI/lqVSxhNDLPP3FkEyoHaahyjN1DWssYCX6LiXMi9K4UBXBQyZvDI0Fo3/NKGVDUvsY
Eo3vKWiyqBANvdOB9MpOnoB8Wou5AYdHEK8CE/FAar6xEYof9GWvaMCIo0iRay2FOpZWhvL5Vmgd
DkrVDTcoDvesPcxHV5TEpE8pI+M7gDr1tOXO18ObFNLJ9Vw7Mg/qjzp4MUNEwxinwd97Ao9a7mes
bLf8z94QO+6xKyADM5sD1nA+Yh2jnxXA9c5oyr5/cq2jViaV3/WsaB4M+qKhRHllrbDzbNbs6448
WBjdyvnStLV34xpv060MYymo0iEscoRo5mdfKshxRuBSfBQju1uMdFCxymeRWMcmXdjmkE3aXkLD
+YBGw2s2/ysU+PDdjE3AIffdHAsnzaLqzskfBpXTP1eQ1fcTiHyMMlh1Uy+gRISbYAIQqj0q3tce
yXuxRJ+PSea4jajTDFc+1fBDDLESyz14WCgVByftNox5BmInKH/GDQmxNIS8sICEBFpYckVYKc6J
SWiX2yuxgqcJVcpV91QpfsASZHVgNmQQnR/QWYB8uucN0g+nviQGGX4eeTcFK03V3Wo1GZW1Zh5u
gpAmNXkMSQXxmWblEIYThod1YquZy5IB4lFmaHsQYW/PX7MaW7v7bdJ7xuWYLlIN/GiSIOngOPJa
gHcWiZjA6eJmNnMFYdGlKHiTBpKSHbJGuzZjcX4x1ZIpnOHofwaQNM5DR4St9Ymo+QWKgFv+H/AL
k6tQNSxs0vI+8gIJNZaJtQkDxjoKoNE11meN7ePIQqeXNceaRApOcQirMkAb5pSoauuUf381d6kb
F5Gy9b73uY5V6GYeJmTSYEF9ng5rFXNtquU0I4dF77y8Z21YgwrKBGC/CPGGyABY2ZrsSt2W1YeE
NEFVaD3osnjSAMmXVdQGxK3Zw5zNsyoISYtDgE8G9tSl1Q1sn5QzqfAiV1uojTYkRu4SNhYi7PxV
w/mpA+Orp7Mnd781EwWdcp9IC+Ta7hSoDsXBvISBcUWfwUDW+nOwu//qoLRhPJobJBnXAt9wIovI
/cUrkVddIsffmfOEzTD9BeOWw099CDdJ1hfrpA5GL1TGT8+sFZNtZOiI28A4vMJcoQqarrxq63qq
whEImOyX3GBKCoyLXbuJCz3elmjD+DWCgDksoQcFcxP+q3NTAuDumgUyXb5ItCt0Mgu60Ko1D6b5
mFjPsxD73/lvlcJVTIaR/YilcEzRQJbF6b0bk9/w7iJ1H3GkK4BJXJ66BtMDBVj1Tk6dWrXlNwlT
ZdUIjls9peVTDmjEic2U2Swz9OWDsSBf2MvmdOBnXM0ihLvkjrJtuJsCci1wci+CYJwNCoyrlNoW
24AbklU9Qdbn8XFo3N3J+FGwH0CK1BB3X6xj19iijMhz3x43cE9dxe7OB15Z3EcCzIenm4O93CXt
0kF/0hBsqk6wrVpo0uWLbJNvRnQzaqMOidfoCtg/0CfxfrQFKB1sbvzLZgg7/r4qoPVCAqU04Wog
m3pxWK3X53LjB9f/qD4S308+t7hP3bNAtHvWXkfgA1P1NSJwRYtNjCxm0Kc1d7TaMAzD/86Lrv2O
3SHK9HS27Z6djXkZ/r9o2c96uYBpywXVB2+FJQuVFalLm4tuu3eE7tl2snAkdxj4+J6E99EciNyt
E8xxjUneTHow5e9dnerQojRvJq8EtDRzkaiDU82YXA9pV+bC3OW6d+FXdzw80M3gXlqPliVTs8tq
/zljY5GXls2KprIKKschnEsnWQaIpi5pZfMLo7VwyM6DPqNa4HhbJXTHx8qA+9BCgUXBrU4LzSWw
YAqz0Bnfv24upKlh6Sco0EhqKDkd5rWRPcj1ijVPVAhpUIeij8JFFHzWBgmLCuEBQ09gGjpkuviD
mDcQPf9dCP6LjZnjnIQV3yMAIThPbmkIPbuJlHXLod3i47ms39fbKjBIf0yOEg+XPbz7IDjl9vmO
XmgQB8W0E7kR+yygRvdLcCdF7o4tRmwuAJnQTcBNoyp5EbvGwMzn+e2ES5Ct9iN5Xj1TzbpCdr60
2lWF5LC6DWmV1TYLbXDr7TtPrmxLOdfh2bnD2Ai0OsvSsFuBjLSFhXo34ZfXlPZovF7RTNWgLjep
7B3IruyOsPYmCHdHve9dM6BkzjQhCblvC4CExYPzK1QoQM6YKqNhv1BcYAtcEIR1i3VT+1e24SNc
Fy38MTgcV/qm3PRcPiaU+/elVnmKV54+ZoG7RaG4eYpnEteXoQYhKWadEqkm3nQdT9qC0kjHrAmN
AbcV9H1+IQ+UeTGJXbcH1jnvloV64mH1lXLJtuRN1MLay2lyztbugcqieWHkwL8LTw+LIJhebf+0
p70ogUgiRua/e9w4TWDsbym8FC99RXpNLWu6/mcL25fEkMoY6nY3SGBTee18VycWaAFrsyvmIuOr
2tn1SvBzHo77aFU4aINSBxQkbh9mYu3omi4GHxrRq/dc7hNC8napglLJXsrVXuUFwp3Pnc0oQswD
Y1qLPArDPJReHoofQ19+xMM92bjKz/JH5z06M7ScOCrVuBJaQnujdxSMUSGQDpeSywhqmRS+Bwx9
T8oXNG1eISBlfbN3qZ969o+mKloYSByevKtoWhPMJS0fCOCdUp87XKIHhoGTM/qqFStruS5ZY+q5
Qi055uqO/SEuw3s6DYyiJ4pHzxmMzPx7HtbLspxESeSpY2jHelgSDk8hWpnX3Lyxx4uOwvRLeeQK
AJf3pYaiG9ytY/4ILKx9eg44Hyl3NG1mpDr9dyUnCEhhTBg2pFPf0DUiRkvlquYdR8EnPyU4ufzQ
/XnRkQJU78DEUJ3MNMQFPl//gfJhMDaCntmL2hNJidTdXDyncPNMyvMe8W4ZkRq9S0apWxcgcPrt
+PVZxx1/x19l96kEfCkGchgo9JUdoShwWg2oa1eeGUzNNQL9geIAvtMdlRAnXV87AYw3U3cmeWHC
DvNVRlwK/4PLWWH+nWl3whiyCOQNMAzm5IrYEuy+i7zXtex/UzUWla+znQNQEN3DG8q4wKrDUvyx
uy8g+O4D2xzTmC7i//wO+mgw3+IzbHAhx/RGRGB+X513SeO6DrvAqswwfABpo6ssvCjtnezpVFyJ
ZRt2TTdadKu2IsxqLaol3tkeZBXGYQrs3pWqjapIIeYPZzhpSNLw3SrzxvoixZNAgZMh8JnNOawU
JlC7Q+gKkxB+7jJdei/u3HVYjq9bkUdX9n2zJJp+ZL2n/wNXVHUMA6al0T7/p3YyPh8JAqU8DKHq
2k8Ou7vDuFVqASHyDa1XctgNyDstnpvzEPozMBNG4inuii6y0FL6Ds9VwXf3X1QyNaDoiDBlt2Fb
UblRC0TTu7jR48ddPopZZ4DYjPR4iQrxsOpd62lHt2De3xrBftJLRIVnQSWmGvOK+QefW8scgJj7
Nsx5CVnRnm3NrqhLuVJ8csjX0EI+EsGAvu32rQq0RiBNElb+nyyASE5Z28vKkpPHsF0A4GI2hRKI
mm440F4XUmwv7+YGNz66n1rXpeZOjlMCu2VmbIm7/cWO7J69DWAa2FHnGVCv+lfhZS61d9VcJSQw
pJbI/tcA2YdyT6RJKZ3KhGBGSpE7KNA+L+rUQWy4621V9bnXQ/ftzH29absbhySz+eadVtypTqiB
UvCieoo5OUTFIqqFFoF8nhUjTDnAfBfqGot1kzDAX9tmmAfVgeUmx6UU5Eew11wz0KGIAki9bonI
02nea9FvT887M2/HfegplwpaBat76KOccr3Zd41S7OVt7X5pjAFBUDgjJyxqT46kkiBPjBIaA3wg
O7dMQo8raVebaRBR2EQVTYjpDjuV+GD13hvDVDsaQUFzozptGF7BFiW31YVJOzfWwUNnEnJA1iIA
RmHy4++/voecUNq7REdhbe1Z6wSdUnHQVOBwsV5ebIeDHOhPjtAbnEDkpqCatfDKthJLPq7Ncq2U
IxPmgY2ILTXN2wtgwmXDsoT5hTCJ9ipEVALjG2JARMBl9m4QcuCLt9k+ZlIfZ33Jd00ULPsmYBsb
a7di7kNhVs8nc9aOfPd/ljsLnRE1UXQJ/vvH+w+JpujILcrUIR2sr4HmpoacOQplcTPw9Kyt7p8S
ZdkbzmEmSoHT5OBfdxegKrYwzWQC1l8DxTrIAi2gy+DgLbplZo90jEuvgXzOzBJFsCWk0ir+nKd8
uaEoGHiCPilLGlgfnyiQAh8F6rc9ThS6JJEwjPyhwU5fchg7sbnQ/Ja3KUBaqeSVdJqtP/ZYB6aT
1bqjZXEIP8kgGdAZR/L5+jWGNENGicTAwR4EI6BBDsg9hQFlMW6LgR8bRtH/VyTLmcORCi23QVuq
dSKRReNvNxEQen8x7+bUocMnuVjNUEWMEshzkhnBsvnmfE33H3T6cjDz2g6as7nBi7u8r5yflVOm
MtJbGv/kQH3YNb0/axiQPjgrrqOlCMsD1vOtR4ymMd3Tw7vWr5BKfeeaUKaFNdW/q2ImYnlZijGW
lzOJrYa/RkieJyZzExyJbYdWwK7ONk4kndBsSmdT0Z3IddFXY5FLx8yq4COKSr62UvlbF6EVGKeR
fpre8/7gMzSCoa1/ukmcUQ5xnDSBc0bfeUynQ2a3UcCXR6C2QiHVNiOJt1gpZALEUWs/KjSqHahe
rWs5UK/qaE2jPNtrT0PWOHhfmLygo/TAlRH4s6KVEbzgqxEKZfTjIqE0Y/gHeW01q4+xL5Ew36Ws
NUFQHhX0fD3ENwGgBqZH4p0ZUd7fV0UCzgOBkn5ZrvPbcl87KxMKAzvdYLyjAb7XfigUkIcm90a9
Cqi4BWvoiOTDgYJKrjT0i6pZ77EXOiTlQBsDZkLGDEq8/vBXKCqrelVQXA9y6MwthMHXGeTZ/TRT
iw4G46JG5k69/vehVaP04CHF38qxPCa9aQj06fm0tUN+IaCXO/Je0Nh0P06lxznZW8IxxcKrmJIo
PPDz5z+L7BHBU8p92N6TN0YMPlPbua9GZwC12sOj+M7a0OmKtI0FT15c14UJzqRfHkX+Dip+DO/5
jbIQOHKRVc+wXuftzifGVUyAR+zgHSzfOLV/69WrhSfLj0ARsRGa+RVmfAaW6znRVUrKhEv3Jaj6
eu7fmBDpcaQ1+tOrAKSs8bcqVp5ca68JiYy0bOI+2ZeH65gtwakj7jyTxPjCTyxKnAshiefAg8H3
T5kNF4Tuy7VT1Yjcq/Axw+25TCCq6dREJtxqzhP0bJ2+AuXIA4qlTnTXx0kBj1Rt9ZYw4Zf/Bgk4
ey3W2ullGT5UuKdKb6Dj8uO8gLxFgUjTQGg1eZ5SHClBNpAQudM4mOiT0Da6Jitp80DVxdnI/zQS
Hdaaqu+yN0IpdfgxxlT+2DePjLtuW8dOLmvYCdpBfDgnDQGxbf5QwDROigeV+k4FY7mVqGGBTDee
GVHRdH85+yw/ortm/01sz1rAdO0f0cL0sor/xEg+HER9yl4rOUC3qS3G6ZvHjtSx1V9iEUPYS041
3ZpKnZqxhQno/JxiOmuzubjqX8+3BOZn1qithZx86hsKjfm/zJeupcZxP5bpSfwsthBXT4Xi3oUE
sBW3p7b+Ayv5Y88DT2P6/tGiNxLJxfZIyDpGglQlQ5klxjjn7DmNQJ1UdvoovuIJp4Qx+iF03ZRX
FwlQfzybGV8qez8GuzvhjYTZuykfAVFX1vT1MbOd+FcirIAmI8EXGyHisgONnvlwMnjHcltmqcUt
Nk2PitunBm1aUFjsAHckpAFuEWUlQ/8c4nERWfNejKUp3DQ47jxzk/Gv5d7S5MwEfhYwIUz3BSDE
bMWaonMw2BlnbsSM0MmCA9ZXJ/FzGiqvT9A1civ7LW5ULw5YpvFdlYo5bbXGA33+0fVIVu9r7ZtF
6H0KgSeucxDiCivv2eeTySZos1TEzXzAVRFZtySO7q5ojVbf0EezJG2iYM3VV7qLpN8uL8+9pAA7
gGf4ObCTFqpMeShcafoM9byclEN/EA10l+aNS9QuIiSg0rpez5ibyg9tdTzESgW0hXxa7lQaywNd
6Fv1csg4V04XMG3Jl5xa/VfWQUVuCsMbfmK33dPChVvjemst18BPakI+gwneL+v+Omw0tSDHV4cG
VxbM8cL+/7u+8x/SjktzupeDrqqIjpJXg2svVVEAJlnDvWtaKCkS5QuEgNvT9+U5c4FkB9C87LGA
F8/IE+4JbVzEXGMglAAuoUw/avZ/RTNkuJVQvcDbhEyCcBoeG+FyLbdYPoyYEZpBVaOzqIM/7sQ7
tuj60t0O4wDGv/J8QAsY332kxRxxNViwlWTT6hPsrusAcw1TrUKX1xbs9BsBBoEHpqimlS+Bl9zZ
5WcQ1IO62CPt9tw1BIr1DHZzyaH41HSQzzSR4tkRYGhYP6PJT1bbo76aaNa3DPNkcZV1LEDBWId5
hmlqMDEfh9Dz3vwNs1eIvvKd8mfBqfbtHqphv2Mgr3EPlQObP7h0pTul38J1Ib54ICiabY3FouBF
og+N9b+h6+4f0xvMF1HpeEfz3VnQaHnxPZ1H66zzKw3HhmabpOiRzYrPHP8M+H4swO1ixz1OeKny
PmhtJr/3sSzcRhp9GPELeYDh7To7uUGS2AUAgycgmZ1S3jk7ZWRSQ3sQ+G6eQDAE0Ak851y4h6uX
9ZF/qAyUreKwextujYjvd3c5rZTP8ZpzfFdYscwrP+P9YDhEFJlZLeFcrCitfEU1MeLpgQDHWHAw
0crcSPUzw64VoPQyuO8gOTx+0eV7ulyrlqg7ikQOfrbK646qTDe/zBK+qzJgMxhMlE07IS+tmIz9
0WDuKRgsSTpiQAP45l840ZAHPOhkA+U7p5bvja9NA1wkUGn3lyW6f9mokBle1E4vcalxmBpjE2zO
Ai4lDvrKjKW1aO5RlCMugupDBuctnR1sKcGxEwim+/+2OikO431XYAP9baMbBV1mFv4+yco0peq5
cedbj//NlkaaPwPNLsVi89mkHCpXWCsKOGro/biBrfmfnXJ3vT9i7kjyQm+ZsL1RPOMp8rMMlIqM
rGQ4sCsqR6/UWR93cZ/yROXz1wMozY8T7SmB9U6a5TjIbfDsIoZJZqPs9Y5RWykCsxDeHH97+ZSD
XARrofz6N1wqCzBaub0P2J7HsHMqbDqGi9Rc9YiV698GnyXjwe6tLJ8fdWG392Tfe9+eZuUldrlY
3dlDKGW8p8j/sV6IXhnOI2BUJDUZeLoFanlHYwkxpFCw5Sp9oSvy4x50g1udRTUSlbR4seWL3f86
zB+HpAEAI7sQVNnpQTjVSeK2Q+RxPzCYMLPB5U0OCRUmeu3yvMBOoyE1M7Ki/SIukvzP9qQgGNWg
uWVRdYcBDu3knauBH2ZCn2yMCQY4uz0M10AJtysA3yA1wVAT9/lo6cEuiDkJGkCEhTAsJbSKAZ0E
xaqNjatF2DLEh/Wtaw2xi1hANoJKqrhuCnd4qa0KKKPiimWjlzkbeHmtFJXyQLVXHWl66HB2oYk7
UG4jDvA7xYX6EuzQqX8pV7qPsqn2wisePeN41uJ+1fCvh8RnueO7LfgKXk/PHFntufY/MSqWGEHV
BXIsh5wEu4gd2BvO18Cxb3bAAgY/9KY1Q6tUqyt5yIV4dF1qouLoj+Ck6NbnAEQI5ngRm4EsEekn
OLULg7NOqLzguSwerqAsbRVBicuDOE3H/h7cyZPKpR4gT3zLYx6B32AxGBjNwPpbl+cSImwiM7et
j5txB7Fm/x+sFN15IS0PsnewTfSTOwrGJqyaBlK44/YllXTljOvMPQDGyZW0tvh3rzzWF4DrUiOK
kcuLl4uzUUTzt7LHJId4l5DdljNrNbDBRMWLHqCKy7oUrIm57h3Q27xOet4pLTVc8tGDCRb+LBIh
sJsS8UZHkI8cyiPM6COXrutBSEWdb4RlMu9hZTy5Zgma0gCK/sc7HrKBinX2rLPdnBZqAtZCi2fz
8OwySs4w0JQfSIIf0fSVEv6MTrdi7pRHMkJxM5r8I291djuUlzypmzq4KbWvKhE0tny/F10ikg5T
R1MBIUb0eXr0ljwAgXeTOZ1bO8V1jND3YQ/xK/BRaLtdteuZprq7+3G+H3YcNcrS2vA6SKnS1zVt
mL1By3vmECzBn773l+CUxe0n1hZB8xfN2DQcwsNsejzfcA7oQ9FHeHUpab7VHCi2rsNwx+poBHri
LWEc70ZEhgLYR4Jdj65EG5rPnyOQY2m9AeTwTTWoScPcEiokC2gW8faMx9/UXHIHUq/ZqiRiryMp
4sv9IM4i+7LUVig6SjqH7F1MS1GSZSTeBNIPzmCTW027gU+/YuaFT2m6efh46QjbBD0CxnK2DD6B
cQhsMx0eTsM2XzYkqMOAAxU3tpQP/wPAS/hRQIMtlDnnyVsTw0KcXZuAQvyMBbkUaHqHXS+845il
kvTl5ueqQph7WM2Yl2ekOg54j61vQ6/yHuaJfKBIjk6pNiGUsyyUqRW5GsYGDQe6f2Q4Dy3Gv7Nw
AntyZO9U/YN5uNRqy6/UNdZoVyXTNFdTsCZDIz5uUwwkvJKa3fn2NtxtVILQ/KGMuYi5RkqKOW9m
2pbuSn+tYE36UMjY8BeRBr83ad1uVSwyMz854TBRXfp3TNYMh+4Y/g9Kpnxgnb/o0mMcrf0Q7s4m
6iU7x6EkMmIJCzW/5vIXS59fxqOjPrGQcT3P1tk+8jVepY+iW6q7JPixa3PO4ZeZO6ywSX9z/3DC
3Iq/VE7PHa7/NTVv/nFjF8BdZwgEm8afPiW/svVR2BFG2rmXNrCYMAvkGagcKaqP2eQMAi0V4bgR
KqL7Z6QPv2IEFwZJqegQNrfBZjBA8FrvtULvNoMPqtdQu/iANEO9mEMo/uGit/342lCMDbDxqkOw
Ji8/d0wIV532gNwt6jfuZVynof5N9Dac2zqfUWwr3evkbwkvR0B8HTdabnIfZj+Iq+50wRfdPF8f
wwKR1hgj7Kqyizk7GMVS69O5riO80TACeBEW0T+v5kGKgMmOB2Sw0fm4XW989PvaZUSf1KDU8rCQ
u5y9Cd0+GR7H0bZoxDdsK07+alum3TP4nIelxRy2Cgy928Kvqw1/y3+G/gjFSmBsMGoOwp2aL9+q
O4p/HnDm09oKw7ZCh4eeOIsF+aVRvo+c8VFgNL5XpOOf6kvGm9Ey+dbx4sDonWVOhhnMqz0Yg3Pb
QF36RN1zTBO4UlFT05ikNHlW6Y0QbnlK5S8YHvVWJmTuEFllRRIAz16Ky0e70aoCwgnPsfk+scX8
uNU5T+cZfXdnnm+fnTUe8o2fyBXqWMITnu2YrefSN7OfGnoG3lD8CmH/RA7WS0DCvDeQ5xZzZ1tV
76Hor4TsRmATCV15qxcZhismMhKBzh2QhdVZMJW8HRRXnu+DzI+qxdxx2bcq7X9Ldo9rqHUwFkuY
qqYwaRrcoVPkG+ahhLi6K5SJKzwjPByds9attAz0ObjxEXjySzCj1DXBsZ1N/AJ+/z6grwr3gtFe
bfKT/YCf9/o7aX1M4GNNny8zCiX4XPpCpacyu2y6bZnKtrj3i3e8+bMASA70CqjLAmeGhSoZmL4T
sU4rHUMzu7e8BY+GkzALqMkFTxFj3lQrIILdNrEbDrD68o2369BZqmWequAJ/svwFcWy3pPi+F27
CwUx0EHM0JPe2uvutI5qSop3uFWS+52VhwQ0SNczcGzR/TQcJ4PpH6540eXjrcLuK05cPAcKX8KU
mDwzQIEGzUqXRYBrUWZ/rkCnlHK7zQSuIFBrQsXtAHZxv8Cl4EusQmcuP8wXIH7b96nyvpazQLdX
lTz4hlKGzwbd3/3SPsKS3QqlXM5+GtkPJIQRKe2/mWyqg5rUtBTGCWSk5PJZWyTpSQcw/YKwyPd+
AIhgrd2u5YBSbvdYImBdRdOvsHnpHqsy9XRbQq1ZxfRrW05ME33miBp7pGdjYCDwSfy2fkZ3b44W
ByKsnVljm6MFm4xkcb1MJ2oZZ89502A+6huGyG3Z8Ilq08ejqxyrGs8p1BIg63LyIBmogwX/wj0G
uA9SKtjMrdkVNteyZyikUZbUjYEGXpKdCyPydvfRt5/uaZry8quWKNmXLO8zhNcQ2tcvA2MBVLfa
vQcigCeMbH3bNkWtEQo1+PqPYkLdH8tC/x8glAehs0K0qy0bqqSEORkhkR12FG0S4Y9GzMXq2shP
45q4NPezQH5JDyBPxMlclikg7j5M2eBClnZfBybQZMd0TNbO/+kqQUfU0vewPAiGNCrRcXfHo9wQ
Dqn11hOYb8g2hqYbLWM/rKBtW9NRKQpU7lvDYEV3VrgcWH1v7zrZYKCj8u+bqjmgpojZ2yw4Ak5e
i2RndfB7LQkh+jfxj4A2gynKFXCcC7c+HVxrKY18eY1pwDHD1cRk3SQz+A0oCim9NkindpAmvMjL
w8F1WZmFFW3IKszPNUKAfabB6C1XZEm7OpxylUd/Pqz/fPeb5/gWC+G61JW4wzrnZOXHOvv1KG2R
dDYL3Fb6Jaa4wbQHgbse1eUUVqrfocUEJO+kuC+AA7U/2kADT3Rh2vVeOJE62uNz6ID5XYpdtHNu
AggIfzrzGIQAu1vsiaNuSW12FHdIwXkLsaHPt7qeG2krnF40+6hNVGW0S6Equ38OyfMiuDZtA6JR
tpizyrNHP82j3dgQeE4/GYjSUy3trQdKIIPxUKwUG03blNjY8arS4ph8cVK5euj/DM9y87lc74rZ
bT/GyPVLa95daTx5Jr9dCR/H9WxAasXRZLRU65rB5EmhAwVtL9yYtzLn2zAuHyZYrbv3zbiHeaGW
rV4uqAm6izI4Oa9wiMWSU4dxAwBs4BEpzhqTUWjYsTn9RTpr9W+O7aGe71GNJMb3czFcGZwpkoTC
wbl+HegSJTvLOTkYhksBkUs3ZobFmknPI9GWH3QEwQD884uy9adqbjtnJvVxukA/fp06wK9F3p/4
fzwsik/8rMq1E865BCRS7GHcS4YRII1xSeKenA5rUaPtGq+EaF/YvyZJlLkb7LzRW9LS62MZZaS9
wnsoZ4AJ5AMGIB31Hd3kiJfnBFZa6a37paUi85vAdGQknl9WshgrgCZSIT/OHyELWahe3cZ/69Y7
UEiQ3JHJjXSReFKXbo5k0rSenMuxuuYREknpi5BRbxCS3D6Dp1ghfo5FCENIWeB29j4++gYUKwTs
nQKgDLDJMIxWy1s5wlr8yKIg8YfTBX4yUh7hkYONQFjuNBfztmU4WlMKWZKjZ2ILtHg5f2Z1COaQ
q8IWpBkDWLdHRpQ1FL2AVDnFV5J8nrFOHCjIYRn0+l661koBezSYylw5cdA5MO0+wHZuiANj9cnP
pgjQ0cXO/n2Ty6InyBopxyxroCtlKF3nJipTQMIAhCImt4QX3Uw6ZwvpgFGU2BX+/8Kw9Ju8yrsz
um0QgUqoMwFw2ZGYbgQtdVAJPSS9lNlTrdKQWfZZoPicRXRTBez1W00fQs9G+Ia1TNgusk/L8jGM
CDDOpZgiJMxAv19gO2jHH5B48j8WUevTOvEbX8Qece3QmOUC714M/uFzHajEvucjkIrKJPEatTXm
XFkKW5o94ndF/+y2X+lX2Ckd58zpPtKmHfJz1QWW/oh7IG1xZWSsMIfUMFMZ/Frx2Etg3vDU3ZTN
Be7yB33Uhl6Fy+ameAMH3W4gLh+O51uCUSJSltp+2X6vSw03cqJ7q/DuEli4l4XEWSSzGLtQx/YB
H5rwtXUJKBjYataU475itR8m4qa9Du0ItWol+TF0KFBI8zdBsvNFzZY3dOihBHxb8ygxJzYTF7pd
obYJ2NXFOO1RNbYEKMP0nsLQT5a7Wg0yFEtZ4uUlDj6GNRNCkEsTCfYVglZLRRfebBHZw/A31teZ
1/TTf1/9KFwyyoqOAqgt8ciTDpf9txhf3dt6K2jiINhdEY1rw5Y0kcXuSssbLwPBfd8qglwxkT12
a4H0VWIgoDE1z05RxhHjknlQi73aKVllXw6Ft8O9iFdo9t+scWmK4nBCL3Qnmxk53vOWj8PE3CZT
p5h6WJi1qv895QPB3u7oZeJ3MSwIFZuDdxn8eUUzNb8s3JfrzThx6idceord+8yL/zMhsZMYUUMo
IKhi/mBJE7SvTiImRvmbAKOy/ZoVx0SxhWgelBh2HSnZHXQzFS9nMkF7LTvl3a0aoxbpxIGWdVCK
Sygjdwdr2HJ8eRZuT89urTUM6paVtaiRddNLqXdCl5kJC/bUzWG3cNbi4A2OHdMyajDuV4YeWPRy
lDUl1gvGbA/miTxFp5NrW/T2+ttKxEJVztBjEBXZdfKTPDsSWPQCP/XFcbs9jyWtS2fmURZjCbjG
AALZ8QfdO52xeQs9YXUnP9EGe139kcQJkXnLZ+VG9cBFjeYm4Xm41AstdgkZUa77AHwIFVCAb+84
c0ormvkg/RboAovQvMtkAbH3LH1veKCJTL1Gmd+GVtzaEs5Wg34nC+w2xDae+Sc5zNVZb+doJASL
sscTdpmpyLaus/B+WbmRn4OO/Fx/rpkQAtTJTi71heqdw7xZJFvn6j2CRHe7mfZWNKgjG8Iljt1w
uMZfL2yOUTSCluw7zFDEoST3pQQlmfk/nfhs1pjdTdAjiIQpdvFySW9zvU2atcG035H43vacE1z+
CHA1pn4rpcharAPHZq1BomVCnWap0pUsmQDfFWMczoBISJIaEPLv69lEP/UWPmO3mcCD8N4RIDfn
6cEFcm5PZzR8vT3r/OQsugbYneunw32dM5ZeIocPOJxSP8RrC0t2ov82cJFhjp0jtS4YEfW28Qs3
d2XKUub6V7BSZR4EGaxwjs/gh7IXkFtalRSs8k21o371C+SwnEc7G11gKZ1YyHdvDW2xfeiMM2Oa
7dHcx0IZlL9H8n9+1arG5kPYCiR84WCIX3sVuGtoSKPPL2VhDsIz+V56UZL/fEuhtHaTS4N4r3ds
Feo3jO0Dl6Kh0kGIx5HLvgvdLES5rU/EwpSn05LDtjmQVFItyj5hMUdRZTvH6ZRhwN3UoKfzvXLz
gocc6EsebeFrI3b1y5Kz3uOaEhEiryPAjGrdmQWLNxVDwu7e7UarEkysp8Q5YKWZBr2FLer43S0X
u3558ScitsRBvCmcj+w+RJabMarxkVlLpnjw5pDS3WSK0kvg2/xoqn/3SoBmiNm5ep+1/wjq3YH3
mr3CAdGtE6qxGIlgStcCI0x4Sp++iNUyC7lPHBhUyIarRxRRg1jgCTesFdFYkOPUOXf1OQe7H/Rl
0N7VUmfPDHk5E9aZ86hhrneCNszd4bS4A/xPp9kJkVVXpFFhAvsXXt2TCmQdniSefOR4mQfrvGK8
fVBgzDlduYRBx+mP+irLrFtTLX3LZVycJdiT+iV/yjp9DABYgGZWR/orpBCN1CZefN14vEONoyWz
2a80bY9U6DwT9h/K/Q4ltV0t9X+Q7BoJk7povTf5vr+8rjrGwEM7c1QFDsDovEeQWYoc5bAc+QcG
P29vQD+kreumiIjqYgz1Z5k7hxmTl/PtWgg/o9ZJWv1Ibn+lz1wb6x+YgHzDFak/HPZ8L19/ydnU
mCibj1ZIEG3/OhbopjblLsx8EgHWZNY9zeGxfq2vrqxvIWgej1xs+cVTZLdiXH7TJG8+ghfhg9v1
SHHcGJyHaRHEA0FEYi/TIRzm0Hg+MmLuBvTxMPzp9oYqPR9UZ6tw1KEuLlUGzVEi8SND1DOXxDKM
ojHXQRdzMo++ix/V2EPijoweOzt8+7EVcvJtG/eqHiPf3ZT0Jhq3ftOzm4v4Uy2dxC49vynm4+x8
P9C+71AxMTI4+t6RAPUAboqQoe47VHGn9Ox43kwlaMQke4mWHlaIfzJj50GITUtfv96TvfJbjgBC
/YUaPFqL1PNjVW4H1drPaI/GRyEXDSQZAjI2Z+DwBw+ZC484nM1vkJmAby6mJNoloQKB/3gk/0cm
ahzWJ+MZzdm8pdUjRIz+FG9s/UlVziI+c3uu2RvP4nwVs3aJb1urJpJmpOB6Cg77mgZT8zAwlGhc
l01xNdUcWLcdBzxBQeuWAJV/4Ad8L+MC2UhtsirFrUSbCNzaphPVCIuWI5WlGOK0UA2q8ffHrC/m
C5knE2d/TnJ6lte1fgDnQshu5HZbI2azRbnzhiI/4zA0LP5igdSqW4uGxdnVRq5tpUSl8fP3VUxf
UjP8AWrt1CPPtnt80ZnbYLV9QsD3UHWeeIZ+L3mY/SZp8WBi9bdRzBczADcYz8LeiovPgz0hvOuQ
6D1hz7zrIv+hbPOx4XwIHiFo9mOA60B7t4Vt2d0sylYJim3pOm4kObG47Pjf9Rs8rLzBvkWPGCOh
n1aiuKG+rl0BceVnssaHRJgtMLShZWZjgw3ijjr6ohiEdsbuqWWDmGb6v9IV4MJ6bqyYwMe9Yya+
PJ5P3TjtI/PALaNDyYvld+aMefraiJxLksP/zPrWSQJ9QAAjPR2s37AQEQQpZOHsat6slBqI/ANt
enhlnbAYTSVEC/q/wi6n5hh3EYIwnFME2LAZ2FNzfD6bFdAKin28TCuqkcSAj2tpejT9za+U+TKt
MGSJhBuUy9iZDwbqJSe6y8oXbmvrJdQ+Ja/3ID5Pl+/bunuWY5A1CyIe3J/LRwPLHwUsw7BXvRNX
YZHrmTJXNYir8WHwn9nn/nGkAGtM56Cbvn2pE7lOkytqwKK9U39UgsI3BufK1AA5EGVV7JD+Yc0r
VR4/2sse8l3ylx52bp/vlcHNBdPS/xnyG6sigeaRg2fJj93i3IIBZwAOvQTF5WFW6641RZZBdNxn
WadKfrVKKNTVsSJ1amxb3iCrNH/HKjX2TNaaxrc3ROf/Bz1Dfhgpnr5G8IsPez2hHTD/k/lcflGf
3/LyFqVlhHREDKh9Nydy+LmXtNqNqEQpKhNKU7Jcr52CfHg/NE0eowDt+9E/rBcTUkSTvJXZ2v9H
IMvyuc8RYWlnDlAlYG2oRRdmXs3i7jOJIqz7cxCWwb6i7xim5XjSVAeahGTAdtkFynTxcwQR6GVP
MfpDdiIvN0cefzR7uLQ4n79ek4xrb/W/gttOC3Nml5oCg/zSxRJBJW2ekDhrcVX0B8KDRrhNCPxl
IuRstGiiB7Q9vRjRDVzGpRLbDDHoRRPmjIGWvT39QWq1NdqqKbD9galiPzZ+m59FgCj9cTtW1Tms
IaDttlqq+SkVftEaOTRILWt15+a+TNwPVJw5JpuEwqVXNJTc0t/IHJg56gu9aCw/UJ5Dlu3/UhdI
LfT4+h6f3IlQ7HFKV6YWurKmKDuwogLgknBNO34TFXYeIx07a9N9XfPER2HfKGYp//puwk9qmCf7
gT1cCWrxwbr/OCh51UhTT7xk8SRgYEZlreelqG3XQgcPFY1SSJfuawXQWN09+pcNqgHaFfuH1j7x
mfGBzXS50wEs3PcZeDBaiQWxoLqaqUmDBi+cbixc7oj6lyVaf6Ft4MmmH92FgDLiwB0bPqiGZLLI
4RiU0BYLYDEzannEDp9VBoV0FVwbe34UR++wYKWfgz5N81/rYFRy0JWuT6rsKCJ63JEKA83Wqvne
dzjoFQj2ld3g/U+xu+hH0YJNP4E0LKoMKg1wtorYCdttkY4lNa2hGyWGOIHmbL/IIAaF7wuZ9cig
d2u/582svWI/H8S5S8JAc9Gab9lHpwdKA/UU6NWjeQ0AhXB20HhFbjiqpB5jtEswfkZLJ66YnuGa
y/wGESBtNbwvdqWGZMJAJuXQt5dwMu7JjnT5l+g8rANSc0m+ZwHjrk0vRSeMliHMWhL5VA0yyrwt
lATgWx2OFG+T4jnootZFafBz7mYyd6EGqrAGOj4g97QHUkmrUHfWuqMqTUEBbi3tGkbquOVq9kxJ
TylEP+8g4s0/5aAuZi/Yi+TaMK4CmwD40+o9zUy0jGpPx8UmU4R7a9S1s5yzWBSnLTfZZaEi1ncR
07Wgi6RUmScvy2S+NIxm+IsayqL5Np9TYoBtFZooBz2RpJUoweZfLhKzrmte7YAuHZcPh4IaRR3e
fpdDRVBRc26UdOViVPtnkIMdEGyWwoKAUSwzvDywh7kp4jwPYXI9AK/Xma0sXIusUXtAOIFjAEOP
XusTnRF2Sql2ZWd/NQtBpNwvtCDIkEneqZ5ScYkdq133qzFre9KeogSgknoM/8dsU1ZVP8HrJQ6D
DTQ/vHVoK3awCJGpYDL1fyoUL44o1iFKhn2ckBZhmJfc37W6o6HlrzyDkF++SikwvYbb3dPe9rkA
Vegu+bcN1Smge+9KecpwFKbdaq+iieVpPzf1b+7Mu+OKe7uZVenXvnQ2FNbJy898fkVH8W2Z/EnM
tKww/roG21Y/7I8fD5qn8ehnOdtK6wyXTQhESXXwUIfhW9dDgfvP9r6Z69iIDUhRf09Ff87Bj/EZ
umyvbe4/RnRxyVDhjP8ZeVvN6/okpyRBi8Oi8NKquuZqvHZ9cvzrTwJGQrHPs+d+ZuE+PGNvseax
t7bZpbwQVU2Wez0JCv77CFYuJnwe+v36QAezmfG3/lND7Kj6hg+jsrzk7Iobi6AXjCzZOTOMWbQ3
nxXM9xiScaVT23leE6LVCJInGkjIONECZ94I0pJ+3w39a5CK4P9Yw0egVfq3W/V4zRw4pjjNWLgn
w9Y7XeLZfWsfmnahnVi324Xf+crgpRKcl1T9JfgdM64QW5b/wFe78nKbQd+N7XoHqZ06KZIUoSJB
C3yPYCsw/icdNMWFezlTjFoUkbOhJZzqPxs+YhysCUZS39kNEjdm92qgw8rLFtKAOkJWgVOxsNmz
yXcn8y/GuFZIqy9sHQIhEXGcghZUeqtn4Zy2ZVVt1d26UkNUJj2OqZY8ds+YbVoalOyjMnMXHn7s
80ja1uwN6cMZtD09J/szUVDE17Z8R6A9OgA9NqHPNePEdfmsDKaAFHOuc+gZBgbhAYgm+NOrm35j
gs7ND+wXrTpwh2Yqph4UzFMWU8X2BFlgeirLh5mCGuQk9avDFM0Bdc53ZXODW8EedczDEugVSCxe
NnYlx7BQyy1wY7WmIS5+gIeHM28Fq4iUHi1TeddZhxdkGmAsmvslZJ8cK/S1JLDybqCrtyjtSpsn
fDEv9l1r4mq0qm9LIwVe7Nm00+5OHZGmH9gDzuAoCfCk5WTYU5IKEF1M/zq5BFvzA/z0nmvhSvgV
skuaLbbTsLaQ1oDp/DFHo95LJKrcMLKLmx8IXVALWNrdnzcetFXztAvpgh7lQkai49FU7v1qAKGA
WXUsbB/RQkyTNYIXKZHJJvGLkH1RPUhCrvJL7JPLJFnJJDm/i7wbF5RpHPnE3xWg5RhPbZiVThbU
p/PHnChaFLQ3HXUA9xiEpZ+gf/MxwoW60Q5syS9TlUX9N8R3O8g/RFqrio7a11mq9sL8vO9GT76y
3gn2mhLlfGdmcYGbOHAxsmRKL4JlioNlTio4HQprH+2lXcmkjQgKoVA0DXVMfcTVJzbBdEbwPD+q
4FjdUtkfk0zmH8E7K1LK7DtN0gYVqJbLXeKaPSKR2pwXF/XvjZ56mnVaS32zl3eXuzE29qKeJQ4q
TeLvaLgtJ06V4PRZore8V1PJiYVKoRoyb1rKkPaXoydnvVHxqXp0PREy2wwcqzX0+H38ZHWU+4rh
I1m6f3UrGdg51o4TRN0O1GsJawH/KYfj3ze2+xxpzzLqep0GmCmexpMUZh87DzbnYIrjlDNtAxXu
QHdLn4L8szpYAiYbzuMkzc+RpuFrJDlC+n+qrSsKJ/do/W5KkR9jnIDmVreRQrGmtoEXN5Zr1Npn
OJocftF6gPoPsBRSKXbck74wvO9fy+vB1W03Qpk9hNIx7C0EvA6uCRCj7X6JxwKFedE4VrUxAhK/
VHBs6zVSnp0pxkHz2QeWaUGuJgDXOJqgbaP31dwvk8v4ga/LvKwiCGLVasVdsiLV3u6ATahKzPHZ
6erR25QR1UceK2be+nPQJr8U4DVTsDWrJD5joiiNBytqjDOrZufnFeadlgNwCXTHWrWdpwPMONtp
cuCIWqvMJ/WQMABOT2b9xBxRkcmFLPWRhK2Z++kNpRlheb/pgoh1zVJXPVeJzeGKW9IqW85iiJ8o
tS0JhnnPZuDBmmAAPwnkoS3ZlyFkHpD0f8008FCVH3sJHdgfEYGxby/Qupl/xiiFduZsY/iFa4Ck
OTxALwukA5rAdIbAv+c13Rpj1kVIJJ12xNjrlwFCbwbt24QLoIjtp+n72+tExxIDgdgcVBHKDgdI
SY9XxyHW+z8wMjES+z414KM9gD3n/hjFwACjDRRwaJoyL2C8rKUnT7V70dxwF7lfT7nrPrk3P4dI
td5WkOKtFmC6idS8kue+rnODZczuNXuHRfxd8Q+UQM2+kkSHxnlOxesfaSGESqbdcxGJrwGcMwn5
o5T1l2ChMjSpt+AfLRVW0JuyZCMy5OKMZqIXAbcT7nfKgnvh92Ip0gtvSD8g+nBEl7APP6raGm+R
CayrdvSQFTRs/A9VgC2x9WmEf75ZL3HFFLkSlz8yCgjMnJP+bW9pQcV1X6CBOAGy9OXP3eMoamEB
Virl70YI82+eNKwE/7AQEfJXwrCZpzxjiF+BFP2VeSn3h0diVnX+kOXySsZG79aDQEvHdW6E7HWb
oE5LxNr/co/pTr3QcNJHAnzfvR9DPb3JT4z//yG8KjqOQ3He03uV9EY+6HQrhZTn7R8YzTvHchFf
2FbbHO/nUU/AbXROnHKCvRpjggPFphkYoADjUFDirQoiS5wSuIhJMKJPypwYiT/MwwxfYBgJ97u0
tCNi6MhdonQEVU06uTXmyVsXpYlePAo/Zujs77vvuwq5clirhQ/70c0RPjM3tUHG5KwejAuKu24r
u2oFymGkD7kNZWaWkazJHH1K00dreJYm/1whn7veDT+qPmnaP7PO5+rS2lEq4LDXStPaottUu8IQ
PvxHYM/GGb4mu2KVZAp2pZDuY5DBw09ifCLsxHDOfTMDoTm2SAxxpX1/q7EM5j9ah7N/1uoV/uhf
bfW6LQmaDu7NCFoHcf5j1Uaq+LdFwjW4zCMqSaMjTIgPz+5+GJCHXej/fpV7nSuVxu/VWxiJ4sui
sOqZvtIzl/kivw/FSCzt/dt+y01lcBhdp1HR+xdq0FIce5aNnolTD3SBipik0GBwl9KYM82K/i+R
3R7kBLruoq5sJTZJrkEJQ0WKfz0OStQiwABwl0ISgY3XaGa8pgl0ir/5SKaicd6RR1fkgFQyehmP
EVXVFLaVWzOjrDf2Q5P10767lmrdpcijNoXbIV/9yvRnwuddbxAdKFuOftz+QgbgdyNRg16z+ZS/
T6CgOsdkmC50r+Be0s6s5Xzn1JG71fAAC3bLDjlAQEq/wszKmFAGzeFnP0Am4Y4FNP+UGJKcnpS/
8tRv4OISyR8znG85jyPm3oH4hjF+Xo9082e3vKc4KO1Gc494I12k/VyRCIUb2C/JJpcOTpNYyRw8
4C+PwhmjQVCMMM/cmIlQVg8RxR67UlXGAvG7/51p3KtkiC3DmKJ0EMGN4rcxAvF8Yd2bNz1Pek37
OiiR/S01cFSK5ao1tsWe3mkuASVwjMMkKjY0N9zIxDsMzKi7487o2YRL7kB68SKrrvTXYX+uHnTA
uV1BwvYP4Uy8VtyGaeiXuwOT75yom4vwGqNRlyHpRRNZQSDl+uAjx2VKApIp2dcKTvUksTTmfarb
yiCsNANFXR1mMZzNnlo/33cXlQWNTlepKBPZB9oBUIjg9yRyh6GB6Q5h61d+zgVjkaxfoczdA5n/
2GDWf8l0bIAH9rgz1wRi/lR2SohCmbhN+F9uhWpzHmoXuBXHb53SlJgyp/kFMK7l3YgAdwnWziYP
nh1UsEkqde/tlDzoOB96HefCM0uJWfXjhaKNyTw0uGnxhWPrMNd/KdFNX1sg+4EBbNdXRk2hMSvF
BO/PqAjPZYsblTJph1I5orUFyrkFf2TvxKNyP8W+SfyxGKKGz6bIeHUpR2lKpsjxw5adWzTvLLgt
7arAxSTRFKrulYTiDYKGCG+62qzB39akOBrMJm4bbKjmULz9j0AOsRCjeM55xsuZbckTdvn6xuYt
QIYkdDGl3I0y/6wgMJuvxw2kar7/ejHJk18BuFfa/iY0UYQjG9jxzh4Rk92+tnY9F1g5kIXWJDf1
Ofarm6e9GNtKeO8aXGmdKjYfcBIT8ZsOLzVfFOSqpNqS7ewKFumtJsdUxOI/juPZcKi8nL7HUYoF
AffaVecLiyHxJD1a9tmEFY/TNOu5Uq4uyV2/bpDwXDRFYi99EIpbUeuDNG+iScoRUenuL5/z6UAr
3JWCkuYesPuZfCmbBHOf2SaEdmTd9TDZMyxUYR9XQrT7XxdgRUDFvW/pA+Rq9y7JwcYrncZKnTTH
ePmJsl8fy41IOjpgiCuqG18C7S0fGLhE+10c369mCKfmJhNnSqOHUJr9ghpJJsfQrSh5YR1p149T
uXHPQglkMxK+zqRiBsGSWe0apqZ710GDwUZ3HdJ9hsSQlJbHlglSBpM7ZTFEckpYIW0GwCGyqDh2
dnElxhymKtvBrcMs7D0DhfKHqf4AzeRq/g7nUcYdi/bDt9Z2B1bMqWSB5MzIhhxOr++nDeIdaKSM
idAA7E6fGALNUOzocm5yoVfMxk9otJawpk0iNTJH6Z3hM+R05YeOwjxPNdO9hOVXJJ29JZm+0Jj9
/ZxBgFCVsUkdZG0vXGZLXRi3aMxZEzqN6SYn/RZp8kl+/kIJauVRbcdy+Z6d/G4vJyTy7fgyww4B
OOmd6bDuiRxH+kp1r9CHpUPRzZQabaJ5pTZRUM/t2UkoD1lUU+gkTvZk0eSWkF5kdKBXNrJAGnvQ
+oWOQwPFdCnVUmvDU8toO3bjYj6dSiDwsLYafWh6HtP7pqAK0Ts7YZ26jfkFgPj66rpBCAwMNtRI
hiPe8OzeI4e+FaH9pYBLp2wrW6vISWMOhDoYHD6bgRmrG3jjVqC8KImsOHGKYuXCB03Hco+hV13B
6ukk7FSEJDEnDGcdhJnwJWJRdbEjFf4bH7FgepKV2FhvEOupn9r100/ygSuZxEI0NE0k1TlHAmo7
W+D9NGUYhZTUQpCK9AoYXVpZgQV2lGyANvMy85z5ACRraH5pCbf6gIeqganFOH3nDI46S5L7HTGt
5RK+Zt6Ds+qt99T/LgppMlt9GuTMdzOmyzsGUVBTwpV7oPlpjG1BMBZFnXUGGpfWaa0rZzFFU2cA
rijMHvjar+nAK/zpYD816BpzsP+FbLjiVl9vaivSSvm92GAl2GK6+AOBlWGIpURhyyunigTdazT9
AWvBIe6knxjZEyQFRagyAvmRtSDcFu/j1hEs8PQsQI4OHyDgvJnHjQBZRKDPcQ3OuRHI165H5a/d
FEwHj4K5ymYazra5+ijUumGk9R/Jgi6Svh2a6kagHBJZeY5Kqpq9muN+cqSjyLVWl0yktdIdegzt
jaqSrOWl+YxlsYOUcnPzGknfHevBxYeXnD0g7JugBzZjJhzqBuWBMyAq5zVp4QABg+wFGvExzwzW
ZlOZxnsAGxdSVzOktBR1NBNiyDOU6xeWKsLHfqdEgpe42FE8f8Wf+Sq28Q0cmYfxBMnq68h6NVW9
r5TMudBqVtixI53qe0Yv7czVS6R3aeXxnckc/gIAv08TIsjGHGi7gOlM0LwqrLod2KVrtMGk/hSW
jnw0Tpb5g8cTH8ce1lq0r0DU4c2+s4Py5vDlFFc/FchOyPrQ5YMe7am4H6YIMGa50H7H5Aru6DRf
G9ot26zhbNP4aLemIjJtF1As68DGKM6dZiciGNiNr8PssgqgSS1KnLXrJpn07a2JXEVPic7YxXSh
mvq2591v/vrFwavkf+BgZ7xBcOzFp5kzNnwbXx6u2if8ezAZ8yAZcGbAH5QKGlumvu0ohcQRkUT+
5ffLPzqUgSpqmiNkWVMjFbALD7JngqQQ8UYXlidncJofFOI0p84PaesYwWmNPwfY071ZYplHaF0+
fQgij2P4yb0Hgr25YFNYhA2BOBVnNvNRh5x1WnKhcZugyl+qsbwcY9F+l52aJMptnANEaVb9wfjS
v87v83+eonjcNQPNtL8k8jKw20i8h3AiMNmJKsSeiCDetawjkkYwqDlFRqApk0mpgHlIpVn7GytV
dxFORJ+5R9H/02/4ZbrxEpZ4JQnBW8Y/stsutj2uOrWHZDArRU78eGa9B9gl55Fj4UWGst0N1+9W
0boMyh2Vis+xeVsA9mK3ePmU7pa8a7QIeyybrP7ET4SWYcvApNLkfoyR3rGpdhB16qgtoy/Pv8vH
jymaVCH0qWHCdRvdjfDZE/qrgkLAN3bLLDAbxdVGFaGFIMm0DRtL+E0dU0sWxhj3ocY4zhfgPa6t
xyPgkk8qkOj+nJ/XiyltQU4kDAOppkALSd6BPjMQ9UOuSlH59ajBLh365eKPNyQUAWr3e7K7f1bj
+2JVGLg6jUF/ve42BaNLkoTlU5BVk6J4jLJmmZrrrSQOwQC+t/ENdhUcVbd/ksQdyQXMOWMCF7wU
fsZtBiUbJBSmqedUrE/o2tgsZsR8bruiKgsWt4AZhzG3aCGRR4yvy7Ty8ChUmNhV2tCTvKowEm9K
A6xrLCP0v9y6S2EaOBW0Nfjv7/bM73YjMmp+dJO3wpnIYz8YEoHB4X5K/PqQZv4qTc91UA9LlWRa
kLaDClrlBT+4A3nfX5a+hI5tKbBnAvN5J/GZPIpFQ7VhMgrUuf1IiJeraYgtjwevD5u0r+Ezvr/B
ELDwY2WCQ2pq2ENU8j+Gj1Mm8OShnpJ7lquE273iR4iRuKx9lxgJAHbHgoxz3Y0tXuDz7KPuUdAP
2CovqYf66lHjiO3oVxzCZX9roCO5jY/fioWr3z3s7x1anczwHctAn638Z+QaTOiq1mN8qr7AR3yP
uIB9UBA3KccsOJLlUdWB3gZ+ttoGsd5aILUH3Fb7USw/+MWwE576wtynUf6ycWuu/Blv9TgJAIXT
i5OJZvEmr8MueUhWw0SYbD6s7JazdrFhFioYAQeVl8U1P+7OZ8CFIsubPyauc5R4T9Zo5C+/CBlF
we+jAfVyZAPmS68hvubD9GHoAbUo/7dbyMOPBQCWlu1VNym8H7cwOnoFlMnCGXjPdgwBqVndmhl5
iR1XBodAPgZ05zUsRtKtwPEcFCFMH8kYTGztfaNpzBRQcbZCYTm9th6LSJI2E5P30NenWNx7xrVE
iF9TJJOinWZJlusqu6L+MMSJs3mTWf4B4I75yKe/c1joL/O5MR7pZE8QNpdE5VL1lUcuQf7stFl7
z+dSNpi61Eo3f4Lx+mSEc6tUUcPnvAAZ2yvj2y+1uCnshJGAZfo38NsdLshZI26bGmtnBixX+2LD
2YMk4HR2wT9DpF16w9g5Jg6xd3NUG6LRp79IwYx31muPOxKGAB8ghK8qwGnuJvm7K373ALmsNJT4
7UdSlzCdxpJZI9tI2yR3T0fz1rQfjf2Dc/Ya7X4Fb25viEtdBEJ4VTYjc0QaBhVnJOk05L0phuIt
oaPJBCbUwvbAtjNuOb7QVjg031Q/I1nLrFB2ppm4w21Ple//LmrTyexS0xmFmvIcRsaJEgOYFEkx
w68osHUBTloPMPw0wdI2VM6uWgcf+WYVP66HRB+xZRMBM3Yz5MSHOkQv8r1F+k2L1c9+KKGrQDT9
jrxxHBBRWMOQWakxajW7RaKbc6OMdOx04sWoJ8BRECZIlwkAs3Ul4qK1YAwtjwptjvKm60/ucsMy
b/YyehYNDAET5ivxOYiGZenZ9H79anmCtAXbvIQQm/sxrcbu43qAcYCU8UA3ZPKm6lIHrI0Odm/h
gvh+iNbAHcn95eDWVBFfoRuytq3XRBfeFAN+GW+bUl9swpq479rXXPvhVeP/VF7k1JfMB2C2EtS6
tvcCEsGrjOHuzj0PyP24mA47MBfVy3apzJi1fzwTPg4DmZ0m5cZI9ZGwN2BGMEx1nRB+2dEiWAaY
ud58RBPdBJsye0RPUyRs4cmRnMwVMEyMdLMCN5PkpxGuieGyJddr/OrtAHjzi+6QDUO3OyIU5SE9
l6ZlJpIRSpoBXPwV8F2ee6KIitlnIM8766wDsmEAhgpNMSbfcc6N+WLkN7iG0qdHePK8jrP3N9uu
6pOv9VSQaNOo1UaaivIczutCTTJX3Sa2X4QsggegKTFJKJjcVn5+RJmFWJ/8UQjKItBdEwlTSnoi
avd42/ipVsRfTsl84Vp4fxQl/+OH0eMpUPQ0t6I17R8DLGtM9fCMBWc9SnvZhB3rjLAXWwGK4Pjo
wWeS7XhH3KF/kDxXD4fZysd0wJjZ9+h4QxXtsc033PHHnwNKcDyHDROzmtqxg/SF0+D1VGwWUQlD
YrKVY5JAC9D4AGrYGU8EINGxj38FapClYohPj34qDn/4HEdSFZtQtN914/8DYQUUsJiaZzvXds5u
KujR7QCgZHRtcrijsYdk4iPCF2UKo/0bVSxQwU7H3AEcTPZYkeNam5s9o6nYHHpomeb/huP3PrbY
7pL8LJ3l6+aux3OXLATKoVoYXjXtuOkoDDkmK4aUr5KdVt7tzr6PS3opdC6ukDEp9B82vKCpiLS+
jQU234apLefeAphaS2tdSxz6ODWZ2/qf79ibhrFlxyVY/hJ7I49ch+XhCvabkXJduYmDEJOUbsXb
xrGVBYBIioREdC24uZ/7JzrolmbpkHTqH/nxC4YHZeJGESOm2PAeVHAyjKWU/VwByPC5EVW1DO6x
ovzKUWU/gpVUZs9mo3IJXh70UjK70+b2wUSvyLGsPlAS6495yUzZBndItcAybef7YDr3ZHRB98Ef
JQY7CdmAMxjMlpFI0hVQi6T1/RL9/p5SOtxKUI0FsXpb/jqA+9bc3gI5OIZ/GJz7xGX5i+7boOOw
y5qIGuzYiNv2avIWoRDTdWXocKSxKge0n6/OoIrlYssDb0TYdeoPp+Q09A8RSJaLmrpy67o5uyYw
f5n7JWZeKpbv24axIuvh3+klx7PbsYlPUH2TMrxZWzn2Xq8S4APQzRgUQpDH9vEp1VYPeBMEnJGO
MtQt5goDmqSa4iqIbqXZ9QYG74ssJQv5LfJrKPUvZK1kfuqfrhIOb381dKdpqBWZZHslEQssli3c
Roeo43twYl3mGYb0EIHrBCBAE6sGjNlalfRnAwAZ6Fb3o4z6PwiGYR+KDuYLYTql4m35v+989Owl
dUCDlQMJq00OasttOauf1pSlM2aVW/ubC2f653tu8HTqPyWzH2/W5KKLolXMN1TrilpOwe8LmlKT
ETb8L8jHX8QLnhd8NKsSNxFhT8AwUBu0GcO6VVabiOrh3oD9Y4r6pf4RRd3rKR16M+oSqvmmf1K4
FBcIIMUSAoU6l99V7ufT4YuI9HIh1yq822y1m+I+FIWbVu47vmcpGtBg+O5FFGlCNP4eKBQ0/5O6
Z0LD2YGYobrMPnDw/v7iVBv6n4hDt1nKa8H5HG9qiyyDrOGE+e+MA+9+3d5IbSX0xerv+TTx6VE2
9sfvFseU1/2ShNP3jZBAOTrRXd2ObHlWJKLQ9+o359Txryb/E0z7OgE29LSFjKfNxggDfvDl25xV
cbEZhi2EtB5h/WOFHJiS/L/lDK0i+u2pQTXW9pXG0UZz3+9HorT8H9AXH3y1hFK9tVmbThZZWn3/
mq3hFLvsF2rKeQ+NzN+eG2uDM7tNuZ3sEtzx1Z6HHaNHXADRBTVRemdl8tD2+IhVuN+xd4j54vYK
JRybZ79JlZV0RXHqT1i3oHHjcw9H/d2efXOLhelE0nR4PRPEbESc97qxl28Ck/5oRu/2tCN6yhja
BjHL1aig///m9ehfQxQns3MlwLeKp6Lcu5LNXCgqtfbMuKqJzp0QbeBKpl7Fb38syN3b5otAMzbP
QtgGkAKCWQobETLXoPftSG+abYVdj87mQ2z72aYe7VXK/uIr1NcMQ5INFoAp9stOQ6V3zzIZZeye
8iygMm+cgin4Ktn43RfWAQpb2Y8ie7tXLuVP1LQQO1pdFxtZzUhn6qjbDvKAh9ORNcT3hj8vB6ak
ijfP94+yuO1vri4HUtSxA2qLtSVm0pt5aBXXfcTBD72Ni8DzadKdREKbNtn0dQuKj7vyZuuizcL6
IIHUe3swyL7uIs+Lqz0fEL93XzLY/5nGtdehta/otew7/sCK9MHfE9mBxGplilpvtSjQHn9DGe6Q
XQoA8CkWp7QVfx/RwhoSfarnvMQkQZTCABM7eZ7QfG6wVcfvP5eq/8cdR0Yc9Z+8vLaHv6lR9ilD
TMu2pwFXAuXqD5DzHTN/C029Kza1tIuSIqav3rSSPlKxD0EGn2cHKi5sbVJ8QcPda17h7NZwkVjf
ck3MArM3h5svfiDpO0rvm4IWKfiMOQnq9aHZQi4RiWExtkYLRNeq1GV2iFlN9DkkZk/uRhQKYJm8
d7QFp/LVwqqwyrwQPEhVwgEBmzWdNcbpbllcBbpOrgIHxVrtgQLrCmwF36ftaHzeYcxqGc3EMJMT
ulPjtSEXtiTZE45Z0taQBaqX8zRMk4GdlLsHksIztW5P4yWZBrbuki+lKAJluC+KSz95T7ACd2K2
3pxF12ghX8s/+Rq9TihPpjf00/EIOksOir7hcYeGgmTJJs+v0HmBSUPV05RMXSPOPLnDjY5kbLVY
hPyp0WelO85jWc0tASWP8NBRK/VuIxVFAy25VhiZJOqeQKoUrD7SETLNgjyr0F+Z0Ix3Rxrg/pru
2+siYB4YDsDAhINbZ8hVvUUalxM5sk3l6ar6naAYdLKdQdwJAozM/kbDFQn6ViwggfpiLJuo2HZm
SYlSHFLqpXKHKu23HOghr2L4r8rCDdZ7/3w20iytdzqq6wAqEQsM8MqG+Y/EeDtZrd3dSscACpBh
bZQo8Cyd8VPZXxr09U/4olHqtwCUuZ/0IKXhazXzOFe83C8L+WkJqFuSGMlcKCEoKNI1rj9H69I2
IGHrn/XPCA6xVCaZUMuOBaKGqi3ZtP9hRcr4Tk/PBBwgHgQ+F3XNu1Kt6SwXoLQ1u9zlCXCQEanS
vRKhHhftKibdM7RAb47E4T7N++1/EboxThCeNYjzK9QltnMrIBGJvE//3IJfspKnI0n+sfJCmJtR
T1kJXlgq3qnGm9WXX+NMjpVpFBGNQL2uO9Z1Q3+OISqsrph8jFTG5wuru8bpC928PJIGwQCVLDlp
/1T2Y2ifFZwujKwmaMq+mRl8bxU5rjieHQ5tqvParAy0Fox/Qo8BS8p6am1cBmZVunUcpR41VwWy
myPaFs0qSElz51Q5W/mpnvd7GyiEEihsglc2SycHzq87gDo3s84ElmlvEXZn7Rlu1AmBQedL+gpV
u5Vb0TmE6+C45l5rZ0ZYZ0r9W/wLU6V+4JKssGwhnD87otvkkuxsayQHdwcifSFtC5ELKaEclm+M
jpoU7yCsikgZkmHE9bCj/2rPC+S1dE7Hml6DXkhguf6hfjl9ktMuPBCDdjQDXVzzRXqyWx4OyukY
KCask/TSrvs91MdCHd279ZubnGd0GeqVbDJrvK/SS0ECBLfV+50nEG5sP1vM5i89RlrdNOHtI+hv
s+48SBcr7TafssMsKebi/X77VwxZk+6zD9s1KWn7bVsnm5A964ZLeBOIDM7xFLQjIOHmRAFYePVA
KrqyFK1vwwfXUrHUrl2pcPGBsptDEd/IW8CTI3TfwB5PEWTMRWsEtHztK1YzNoe+xAafr5j1c5MC
EJI04WHZwXEBnICDp4W6SkyyHyk8ZbIzFIBw7fcR6pq0XjbP0FZCLwRyIpCtJkfBvhV199UFiABZ
30L0vBrZcvEizhJpbJx71JgjD9ADnCCU+SSNIwm5kaPiDFEdW9w8sFAyVj9TifyiSriQgJ6RdzrN
chRWgoLzQycp62Ry69q1K/vCfNQgI6xwM4UcKLlDs7wDwNUBSwfywdog4dmMNiyRbXYNT2ug7lHM
z0MX8r6HAwglvnTXOUijecAseeSxUdfaJZNslAblDLrUP8pY8i2RID40OtkXC4/UPHG8jzVu6rCO
vJuGElfZF2bQR872vx2xzYMUOt0qWTgv0aOcTd99yQKu8ndM0CXARt/nHCVCbibildV25xOKwPas
uLwgvbWu4zyhfPkX3v5qkjNnqNlulluJGN8jU7ePjA7tdCwYWX41UuXq1zW9UTO5AFkFFwinNK1V
nJn55yM+rR7lj/p5T6jX67Ddmv4IgFNam/F5lg7hfrEKECSRf+2336FgVQGRpZWi8fd8CfY30nl5
LozDTeruCoMEpupqjzvNzv8nv213b7GvHpaD6CQLJ0tKclun+iNTvmIOFtyh8kntGeB74ZgxNKN7
TRnH9O1NN8ph6mrh5xcCWzoW9RzET19zz5fVMxO+hxIH4DpQskpMxsTphPhQEFpoY/3GTMXd8xyO
pW5bxzAG0v4+RBRs1hOBa7wcbmQpBDsCZvoC7ytnA4V8wSelbpIB1PxxhAmBCjjNFVJAN0cRv5DE
saj8jreUH8g35+wn9xB2JpG2qL/mxYgIGGBTVFvi3VQKf9Gea7ZwkP0QcUryW1xD4dBFqS3oeaws
gFyCAnKxGrGsrIU0s6lwLH0aztRHGyYMwpaj+UGXndNwcsjJ8/O2WUQ/kFXAkxUNGedhfz8FqrtL
UzaS9JcWsPLRram4jT1nEik/z5H/Ofp0iwBLmV1HCvcwGuZbBMGryuheVEQnoyQH1ScW2u5FDTCQ
6hsNSRQGB1IlZEBrCBQAyBl52XW5hD1m7xBBGIm9/bBYai5L1TBazzLg02Np/3HistHLcIavL3CY
uZcSDCXO1R97xKLOPhiuhX2YXTxXHyKleM5JWTxd4YBceO4JSSu/gUCmFaVzcSCwJHKO4Rb4YXR1
zO9eJ+WEgBQiCQl+3B91dD685+LYpy09GGXOuO4pEBitN9TmSbeJPUQErOKIgB3GloN9I9uBJG1G
UtjdCi+S6BMPloZ99BGjR8osW45aZXil3FX4pQfY8byJNTn1I3Qn7/16I32jVmegLW4PTrUvTaGv
XGUbwVU2DUQVhocVDGC++hBDNCFR2ZtZtfSOM3w5KMtbXoKdOsC+Z5wxyFQvKgkVrl2WjtX7aJcD
Flyq7KN5bVrgZ5GvO5LXgwohjYmdlfwaldM0AEsAf9z7evwcxFy9r7IbjRt69dc6eE/2bEBw8Rr/
bo++x7gQlYmYk9v1AYf3dYbOPCzNsB7elU/xfXeg3y1QH2UJbr2IsIoodSPPfXzs8C7pgKVCVfxt
291h5Kf94G64cPFouQ/pUvKiA7idSkMWDVATxAMmQBB+CsGK9bboycX86fSFQqTBBNP76l/bk90e
U2NQ6WiiTK9dmFq2VGtjnQkeY0yaem47YRGzI1jjCxix3cPS9umddRLZjalb/R/zVX5D+xUc2iKf
0+f6jZw7FlPYd5kIdGRiaT9c6PWdC6nzzG3Sy7eHkhxlrGE9jGOpRnHL4K6MdPnJbDTqLA0GhUmk
OAHUEkU5r/at13ZQeKkPODMgS7sAvxZiTkJDSXGk9df44kzvJhT+NoFStFwq4JlH6WmWIMbAm7Xb
NtzkR9CFYi1rUmqeD9PCjJSv8gm/F6hqdVlGIWR9BevEVApdz2RyQDzfFNP1pZ0YMMIRcDdIQOa3
kp2XwFQ9uV04GUD9N32RbKRl4mX/XC9nbTNmTS02z3d2N/57gd+oLshahRnBQqSkWRM2d5eqQfjt
0PbIjjNCXVBE6EfUEk/ILrbSSqfMh6whkufjcQJPqkj4xmHdFtA3uKYSNXAX0HAkHwH59qE6stTu
SDolveTWxgPRV/PAyzNAbGqGF7Co/63wD8604N70ny1+CbvArGLqqeNPvtX09YipzMaOQFnk5J6K
oJ/NlqyqqN6GerCzzgRmI9m6fpaX0tvTdw5/7676Bv3AKZgSdYeATHeajcpU7UZtCUaM5G3elgK4
A2Z+I80nQCMeVvYluSMkFU7gN2FpNya8w/92GlrzjDY9M5ObhyTi6Ge934S47AEG+jUuGtHvAgXj
xOHl/D+LMXCvyZU1ugbQJwKvs6XTkl0nbgqZ39BZJuQTP8XOy+ydzI0KhfRo4+GNSq/6HtM45Sg+
oWOS0o+bZcE4ZCPELEYBcFwABgiXInxQjgOEmd4jIdCFCxXV9ruXmwiH11oDTzjlTCUHF11Il1ZJ
sCmdLizXL2we1dTrmwQtNv9RYdcpP3n7CZ4GOwPiEAh8P9Qw3AYbgzSx3MP3BQGca+mGpkLaZ2Fj
Fcw3Jzs4G84thNBzK8HzGyD+GA7ZpaGA7bY/5bI1uE4Eklk8fRDKWkX0xoI71wqnRVaqCX6HrYgm
1kELAbWjsLJHDSkYsfy24FAgX5DYi3hk2cEGjHVMFGY4TcCRczVrrS5y5fnsacYVuHmjLA22vOXR
5ge7THgnSPEkDJO4tC0YQDnfeeFZPS1JQghPwSm3fihXno2JvZwAzI3Jfirah3RpbMtnvx1/GPg0
g+KHcOr08qEb9lPGsrRrrC1hdqtksVhLlvJiLs/coIqE9mCULWHONbnNQgXAw+sdp9ZvdUepm5PY
wvoBor/q9p37a8le+U3oRXqjMPF8P0jTY0/KV7s8TnAUzdDwtPN9UnH4D5rcn5D3rEkULyXBNlnY
HI2mFMWlT0G3/dmgznGgHBU2imbiAqwwgn4szg+/El74zXpx/xvNeoa87neXVgcMmIfMdPgImDxK
RfwtpMUF4fd+OQgINKdL6ckmqvKR3L9jNkHN6rVNh2Ji6hzsnE66T2NKle5NEuYOwRH96jD3Y6YW
PKy9fpQlmVPVGfVSqd0X5ih6X9aJRCO4F6maWZGsvYqv0cpFt0c3QxS08gyGW4GY6SaIDwyAOwS/
aTzNl+S808872PUc99l6DUpZBuaYbzMYCXe3DLThDHENU4Enmwg5DVsN2Fcb+T8D08RaetqMbnR/
hXkmh1dSbF/Xc/orQUaLPJMcgLei8zq7R/gPTPDEGlNT54bt+5LQTl7B1EsRJA+eVe+okuKGx2VK
VoI4oTjrX0LI7uAw3ddqFyq2h22tXoHscSzKNoj5xdZP8aAGHD8xH0Mfx6yVc/I7ZybYx9e26JhU
Y1BM5nY+nZd9oKmIjM4Ccc3iAzz16HfFzL+JIKk0D2GLOFCzxkyypHgQaXi7x3WPNKXUd841IOV/
tI8+Y0R6Bpw/TrBgx+bKA79uLI280Nb6xmHKC+4i0NAwSkB6b+V92kNeS6bolf2NlCHcEGulxTjO
/N9Ll9lFKlJSmuxPDVwGrcgdVgpwwPpa2QE7nqp3x9MsMBgydEc6iQZH/W7TPAYUuLRbmfnYSZmW
tszio7vhjBJsxhmPz4EvyiWcQaY020GKmUbAPl44jkK2ZQUQYEnFZ/OP5cgWrlwXZwQT+LhL5JEY
aO4BA61W9ECSSUA66ffj8008gFY+knIHxQFrCy8QEqjpTK6A+3+vRf3AJ5WTa8yV4fEIzcVCH5wj
slU1GuAqONQ22AttspvPYvUQyUMP4e+WOMwrYQryvveefm9rMBsad1rcUHq086K02I8dZFc/W8Ib
QM032GKIorDvmo1xSCoo+L29MNkwcClAuAEdLuAVd3RltGM2Lj1HM9DVfqC/R+frhrqtSobjtqdJ
K1gLPyNS+0fNNipfNpxgUuGgesSNuUZ7Rn1UapDSC6qC1yv/SqtOPjy5hbOPHdkoReu5hPlzDrhF
vYGDDaL1SMTYKa2bbY/knjJ09Lb31HExUodW2rcJavGFfPwWrrf4ihcyV20MNDRl/91o/ozz63y5
vJH3RyMTZM4BKsQ/RnsYf8xJPjdWjATiaeJlUhZxvS9vFwf1wRc8miSerMGr6lWNlBRxdAux0l7k
ibA4aYCKJavg1qIYqG8thCpyisecoDVGtQJ74simGfbdjb6lgWuoKfbMWYCg2cTbH9CWmlVRa8af
fLif8D5ncInIZoPxWIxst0Bgz5tJb72in2PI2WzO6BigjuHGts9kWov0kcfpUcFl5v+YsgCQdXI3
zNm1UARSzKv8Zskfw//CxtbeSN9BIl1o9BV8Olb8WVRfLMimxsudPIqdgAxsMb+RW6qrG3ePrkuR
aVYwa2mBzDNX/srd2tRRTHgDv0btlDFWipWjyel9nvr0iiq8PwCJuG7AeFJGmTLl+PWaA+jNxJJY
RP+oukTxFsBr5Wc/mVF0YAUA6dRj3IuxYzVZcE/xFinzmVHhvwPnvA2zeRk0rqufK5JZSjXFdbp3
S2GLZF36zhKa+y6D3Kv0d/soChq06S/NPtEqn1m0LXMBjz7LOZj8IEk+EdJMswbrppIq2VbLRso3
1zPZtfI62LVQ6dm1Jm+ZTmBOuis4tiX1jou0jdSEs4sVIh3/Gr4AyI6w8btAP24CQMM6Li47W2/1
/XIxm8eSlg15gXRMqaCFtEdVUWsCVDPnN8ry6R97x6yVt56vhBe3OkE0GKPnYZ+XzJqBPbfjFDpU
v47S84tXncANXS8cBMQ44560qBTSoK/zFyA/sSJ7+oMopPHhgNoFV9kGgFj8SoC8MXy/bKRAVk9B
+12DoB3ZIIuUpdIPdyNcRyvVa8/M1tlXAwA3oJ1rHKldKRUQYKuGNbNzXqvYEemNSqeiK7h780qE
3RhHq/MOfEg6DD3/o8C2PpfSu39sLqMIIviJ3eCud6v4i83Byp2/NsHuRFBWrp+2V8QUImiHobWT
E5dZz/QMfGWZVcW9SDGmeNPDR49mZPmNdglaSedbhEzPSVneVWPS/IiEAeO+P3wF4VOUd2vJSWq3
0ANazThwTyPFQAZDEja1JCcmTwYMC06YMFB7yTD7g5JrHP3Qs6jnx/UwXVEnsvKXzv23C2wTInVs
6MTcXr41XyAMXocdtvApIZrFhTdV1SoPVvgR3s/N2SeQh1nAR4D9DPUJLr9yblimKQqdsqITUJoQ
4kHWBe6pfiVUeTkz0W6ui1ahsBOq55Oga8ST9vfJPsTyP/U42A57ujMd0TvfsXskF32851Ui0WrC
N43ikevog+3ESV3qZ6Tn8j6HE7qKgGHQ3+fBgWBaZZOrPfhFhJrvbhDGqMn/Oyl/MvJMy77ok2x5
y7Ag7HDCR3LwoNRpdGFfAqPg0oBw4COSawnFZcAGN8k6Ymv+wvQBfnB2eUF5V42LdcjFZ2f81nyX
Vp8gRSDLh/YvLFMHm/sjPAleEH6emJy7i66ly1zHnxfxKUPUQuT4CyJnpwO+e6Ya4S5NlhBZmYjQ
Rb+xrxqCk540G0lqrv3B67TRKTU5BWalMBnnkt8xuHH6Up9yvCN2jezndrKoQHAzG76ko/wSpFbP
leHNbs3VeZOIMloYnu6V0R3D95O/BGtgNDZT3GdwQQmWO/APUUHQEiU7imNdFnSzoJma2qcUyxdm
GHaaXKNUbsEZcREUA2ZLX0KGUwY9qBnkFCZZi3HK4e/0aqYEI2w32TGk0HbyC1wioN+qpcGfBfFg
q7w/BcDajm4LL+FhGThli+bNpvvKwXXrvfa4r3BirQ0e+kYMqAhk1GWkUgLHWT1RAHaS8OjcHUyd
I037iK30YX8eMxnzHPZ2twVFCu4dJH7t5x73hb8+0J9CiDipuKlwEZAI5D27tR8LrauKsXkumk2A
1CG7TWMmBP3beegYyqgNkplVk8ufcFbSbC1rAHwWrhscNbuznscKnf3p2n23vkzG01IjFMsAZb0t
Huq3F1+7f5TdWrc5fWAm5oJkV5axgMjJMd5+iNqteEnNWYDq+12eqiJMt2dtih5XRRIA0r68K/mk
J59GfDuq+9Y89dk5RK/YG4PAwBEcQcOGB6FkocVyUg9Q6QbSsq4GJ8ZJ/3jDKbMAlL8ESd2mAhC1
ATFU/iPJISlaKldhbuAH7p5JRlMisRr6mVuWwUlHPkn7pRfzdoPdRI5qGCrJYJLfigs8BQrZiriE
vpzpkYbrpR7I7xiswb1ivkAk/R8qoCQi5C1ozE4YsajYglTNV+v9JG/wSi5QDUo0Er2clY/vE0es
puaGm5/cmLP20R7LKo6f8zum6UADYNGU8ZUsP0hMMWtDdC9sLFi1H764cmVULWffgFFfAcU1DOrK
lBcLoZ0/jf5TllVKR48kqmX7ioEK5h6cG7HMQzS/Qazu30YAGhA1K3AThhv/4WE9Ib+H4iySmZr/
S+pa6CtR55PRBEvbyrHB82HWeMr9tjPBsBb3wN+pgO/C/pqkS85Qz9w+D1t3nGUjweJp6PxNhxpP
pMNfd7hRm5ooR0x/0gQtNvuoQhkFtZi7lbAik85Bzkz00uyoV6HqfIY6HpZWV5TzMajg9AMS0mjF
5how7QVrkt6NHstcWMXaeRuEGHILVnHfHXGwHnKT8WHQ0+NNpjZC3QJchBv15YVpDDCAVZwElQck
PGTnbUjb5wezKR977OsUSL5hSsLXkzEEgaO3ExZQM3iSYV19lmIRaxW0oHBtwEbb2aBz4QXulqcx
YyxEpHy52R8/jx8OM8J7ZOTWFJM0eVjGoqsakJAwQe8a4baCzTYLYcOe4Y+GCsNu9VU8jWJ8O8Zy
KJ+XmHM84zKixPNabzrqJNpD0lhk4QL88/dRWgTpoujz4t+vItSTy66TBZPoSNr4O8uiivPJKliu
8bZDoqjAOPBLsjQfvmgGIMGQBkq4q7Stqm/yS2QFyYntDfyUAUykAEQzIxONfFeipDQke3NKaROW
Yxwznk2xmmahXFNPWGQrtJI86ixpN/zhcGWZjNT1F73wAuul6YxY7hHUypyONnhtFU9iPzbOidA/
f2nbdrAvNcSgupvp1WkTg87DrgWE53nbIFcqS4gamoPoVqs16QdFiJLkOuRj0/TjEK6ZDBKTNjqF
3XEDgKZNQ3EoYFxv5pQmBMxv60CjCFfR4lB/InUKbDjPAyr6TkCezrb2HTCpeB7y6PwhK/ZqpmRC
Y05hfEhXGlOut+1Pr1hBLfPW3ilGT5C0FL9kt/I14JeCGndarnCn5Dw+wrj8xRr5Kt3y8B8knK1m
ZMN/4K7i3G0V2d98pehHkQzUc5lkPSXM5l1a9jvuI5kLmf282UmCexTVO2JrjAf6qliHu8ABU5Re
ti/lVR8bybsOfb9LWDNStx/L9+8YgNlRcRzlxcCKHDv/70yUBbSoEdreMC2IxpEgPTq827iwwj1p
FXCnUetf7YkaOJ0XDcwWqIvzVZ/3MiBtJqbfLCNV4eC3P6z61fBCJQww4APbTR5fZnDfy2O9vihd
8b1wYIUNKTRgRaYkKpN5IU23L4B9zg+rKy4A9XTxOjLkNlpsP8Xq9rHCpx980hUjCDv0sqNhev0y
fxXehLgwNJZIxsgyZT+THTUjcusibtGe69SYgYb8zoVPczujrPQmpT8Qddt4lgb0qB9YdWHIbKrZ
v/QHyps9MWSBvKrTj/h9oROfbRy0r1zHrnMHuPmvD1tekLtWFeCLve1wO/ySTslpthhQk6iv/oAO
snuxDXcxK0ORWIXLSVGCeLRjkUbkgwS1N1Q9/w/gxj0OVMcnSQ29ejTlPjbDw9+sxjDpy+5x+Oi8
Bd2rMPOiN/ntmQgg65RPdFrbCbQ7QRKiRpvrLP4iYYEhmmxp2PziBByrlkcPS4YRrgDuoGUcM44O
Te/gJYZMO+IH/nyQaOm5YVolrH3/sAfqIUKsB1pS8wiH18Us5nQu1bD0/womYJtuC94oH0o+M9ig
iQGPOPW29VF+uqShSXYtG58PYITKegdl8vK2dBlvOX/9hTkjuuv5LrXn9HC7Sueo91uitGX0ir2d
PAcDuCQrqacQclDykYaWf3QlvcevN8NWYTvcwYMPUiX3h3WakWKWYWV7TL4YQopjZ7cy6WXZBQFe
0gbT09byJgcPiOQHg4l/RbyxVeXmNI4jee9nmxlXHAas2oCSzFgaMlkFJpHIRvf/fSCu7Sxj3scg
DUGF6y5eYxsr3d/e19lLnbHwkqyTAoF1+K/YuOxI5RQogc7U2LgRFTplsOHaRqPqjA1xOTAg/OQa
9n7L4ozQuNHRIPoANeOLqpaO6yNatfh6JdmzogzphYTU0rUN75xbWjTexMxolXVT65+nR1UMTCDn
V0AJUcg9kiOwjxg9ez+CXQi57w9WBOPhxHgTdmkFN6Plo/LtxBEN7EBJXD0OVxUxVJ0yn+pO4yN0
mVKv63XGEAe2iPk/q3xbVYvTsdE/JzqELIcwoous/nDK07JygKZ2Op/ZIBzrGVthrqzcw2clkLas
ukHrhF+TpDpqNlv3a8NqMk/VZB07bB5NUhjXIwaaox3oRH0ThaY1w1/fp2eV6pWoMQLq1pjls0x6
GzQ/0gQFoiem1/jukK2zNV4TFgiPO3TUwGs8MHOJxlSMi8V1u6oPpY5Z8+AojbuJtOToQCJDP9Mp
nF12tA4rdmgZZHFo/9GkmRXxOPHKMcSf4zOwA9WvJugl2S04LkBjnyVJmUUFcCnF0xdoJNji7PkF
8124aDVS5ZL4g2f4NGjhpNfHLVHjNO5m7iq9o5EC7vl2umf15uF3tNfKJmMZYbs4zREEvnvINM9L
3cmACXkywvhnkNF/h97gbMjDVxiOYD4Ka3APXXOiKwMY5MQtAR/EmyJWsa99vESwaqRDlelKxg0P
lJBtPxLhk613H7fMMXl40tAdUKrsHnwBZM1vuxIfl67p4wPArCjkrCoFsLtl8BJ+YXzkpVrCv0SI
KClzcG/Z4oJf8Sk8Kg9UMeKSOP6AGbyuUAxBhpV6mrOKjkgJk9y9yEI+VMRTw4rQy9NOjhVkZXk+
AwyYxGPkMcsnpeavw9uYUGTiROv+EXfKqKBZyjtrTBxh5HTI07FFHjuviGL50xQxxeMeA6dtm1IK
LMgo7adZ2yqT5uyW55ls/zHvQTpf4D1+8fw0OUaUYuf7/nwqWubhwm5hB1L6VbV/uC5oy2iNZFw4
W4Fsdc/kxrlBexxIpXUzh7rj0Gjq/xh90ReGlyJFPQ3hmhY1Imh6QOQfIwzeh6OvdxOcR7XTZGgr
yLbiYglWZizg7ZnO2M93fUeE29by/ULLoGNvvz+ewbeCO6bYJ4NC0MNwenslEk8lcbs8lsUptlPj
s7IbaN46xnUVxRAWab5IB0h8EOBs0OHxbe/ADOw0B6drFXMG4v52vEHPnFWStykZw1d66py1BGgw
ltDKhTgVP45dyS1Ll6xXZXcX/+kY6w1sSD0zXsh+en6AF4FyaA6LcEcaQRZB4YjWmS4pnU4ahJuC
rQ2DLfDLCDZILKswRP3b72J0P+1yyOUDJONoshBYbGCNxXZ8hlg+7C6bGYwLB2g6FUqgdu0QSg61
Edy7+hw60p+1s5eXhXAdh49g2iJYZ3MWZk52Okb7BQzyFIYcxMYNb00P2x7TscXnsXLjVFeBOoQu
lMdarsevSO0eH+W+7jHJmECnmAlFKRt4mb8Df6iqeiBXbgaYGFiUwsRkCFy0w0luLLrgzDVCFMYm
7sUvDHJFAZxzo0IJk/fcprBWGku4683Rcb0q4Y89w+HaxgzVhcsCIXKQfaSdqZHisV3E3BPqKNar
iGbEz4HL3PFIfMHMMmQgKXGaCWrUDDYkGmJnbxsCHKLhCaatckryIupOIzTwrgGhzRjaUAq3hDe7
aEoVVwtzojwsLHO4yGr6uyfM0+/U9qEGTy7/3BuqkBNEfOk67hOLfqwlzUt4u4evU5btJwULiRu4
0jYB0dBwNkbcOnc7jtoTgQYWU9kWULoFyIgvjcjWyjYxfBYIUewRIdMM+b5fsiFLQ2Did8ShdWn3
xi41JnjF3dxDw7VTBfxNK7fyqGM52SgGwVtPsHuO+b4m8vkuKFSDuMQbwVRq4JnQgf5XqG6roXKC
gc+S+DtA8sPPVy0uXWbH6par5uvnL6F5VAwE+9wvWs1wJUTHeJStm5SJWLeL3rWqZsfrofQGlxlR
wnZJpslvhL42OXDPAz4yW+Fcjz6vRoZNqFCw968fYu2jyRfcYAZNuRpzz6FAz4HS2OFFS7S+6qm9
iUHCYNf3LS5zvckjbtJYGYRof342ySYLP5yrO0EkAyiSorXs0fJZ0RQYYaRj5aDQ2qcElKL+iU7I
YKWNhuhe/NbjDovwqwxp+atFsB9GkazQWwOsF37EcJGJdvNYA3bJ+6e01ffRsduubw41GnHvcsqa
Z35XtGRhZLbTGoCpOEk+z87iQmaurPwG1HUfLfujWrQt4RVMJlpEpikFktuFqwKVXyBBtqpFMqI4
ToFLkFDwQGj6S9SNy852RD+g1C9ke2cF/gqVO5fTalEwKEukyhXwJmUykAiH5bY5XYRZwN/R0obP
eipcGGDtqOa45+5gowiFbjOIbIJWzEwxsHbzSaMu4dFDkW94kBraHPo7q+/M1cceMzfkPi+jBefj
76T2E8sMVsxIA1hDSPN7x4Kf0JEF7u4ydyWoUBOHT5BKXRRr1PQsc6SejbQtX6E/hm1ipcB99ltF
efO6tdSogoKNokMa/DMY452/e5w3cJuwClya2Z6n6mPs03FRYNRmDyt6pm5hq0nYk+IYnVyXC/bq
nKTAGLBH5JCLaiVLG9HiAUzKPzMm9NjT3s6FCrKtnTShksf4EL+ekIVZGPyUj5pGk6DBVY23WANd
aqrcrxJUCuwlL3FOMGvWGzIhgz3wTTlkUm9XZ7xnyUeXfyhWQKlp+YQr1cqRaGgWkeiT3YN6YBlD
YUewm7QzL9KaMgdkpVlkKSmX31I6lO0SLBpRW2AEUacSajHzsw6bBrOPsinjwdoSf/shQNZK2Krb
42dswVfqh2L5MlJpIyGjcNFGmUWCnnNs5hP9XZ07iPFlfI7qcmxKSsAYGOYZX0Kk+Sx84E9W9St9
uEJ4nHBD6UZJ7EneOc8SRBQIEkMI4rTH+9cBk1bDGXxtPf6gfrIIkiMiKvvXGRVcBjyc3A0sHoQK
9PlgCuCaAI0jHobJrMQKDA3k2SzLP/+GTLhNdJxKBGXYpRrEuaJ1tdyKFLGvvZzgWHsWv0Oc+2uu
kFxJOw+KAP3BeW+yzqKhQJPiYdoFbOIiFI19YbAGuPZLdvVJj4/eJfBtEq+ufbLiOI0394y4gGe6
JvDsUimLWD+8Jua5l1xXYpK8sQHRaCeN7GI7Fz4qjXAqS8F6kzO7S1znlgKtVOmLuDasvM1+6I9F
F8bo9JFh21TVaYS2fjccS3IPgkVJ4cNfoVYnbbaasb3mYCf63jccqAbtKUnnn+cDQ/2rFfzXlQpX
n1N8bciSXVOVEmGUNn5nxTwT7vsyfHiWktyv4BftkOoyVNslgmjtwO6/h3VCNEGXHuTmewMR95KP
w54f0YB7DKkM4j7RTNIjnWFF4O5QgN845BUNuPDxtPojq4EblYMCd+/yxQ9t4SmpBlxZnTF+8dpw
IqjxsvKBoqeb+cJg+8iFm7LZbSsRblqP/IhAEAp46Uz+vKEuT6TjseW2n7LvVjsKtfBt78h0Y542
WKYjAoSAMtWu2YlkXY0b0F1rvpgohFWdG0HL4oZyjH75nrIFX5HRnWmV2/1u57Z6wJHuKBl1Fi1T
M4bEuIsqsyh3b2Vzkka+vR/pUdflySdSWwNw1iJqLMsjNWKzVlENaG+axEQvezNnKitt77B/ChXz
rAjV63OI/qqiBihSfjvpyqtTLoyXd/WbCUJII2iaatZa4bLh7u3rIuuOICz+AuybAHxJypMAEkkf
YIkdh6xK++RzfxWQEWdNWQpjvf88Me8VD3YFsB0qim+6tSmDWRoFL97nVYVHaCXMiMcMXB5APTrO
XdRRb8TLC308rp1irf82Eka8WUmNK4YRANQVuqLf4X8PglVSLkL1CsRwI/2MLlQ6a5EPmKf1gxsB
LRtmKZN996yRg0nVX50NjD2ei5nXdDt3rDcPepqOGQYTBkYiuUFetPeIcOmW9qV07lOjLDLFzLzu
OqkucSeRzv2+iOEZBJFvTfG1DpbsmKtFsNJlTA4gkS1WKn40i5htKExJMDMObjS+RJBEp61gNmdO
sXLMLdOt9vG8KgyTCFhWHNmUHSgxqGXZSGL2Wo0KQqz9yaSFSuzYIoUMJf6+v/sfS24vxiR3uc2M
n8fOm/OpkhTLZn5TggD41PtDE9gW2gUVvNNnAun5QrskHOFwFzdXtoGbyEluhMNeaXAvYIvvJQCg
GvVyv7aZcrd/MvZcB+LwoCEcBWN/xQnBmUVuZqReQgdmeVVbQIKeXoSmgJ6/dj+K6CxFLWDSzQIH
awNOC14ULxx1LOnLDlrFrkFGIANSReYH/z14wqRq1Ze4lDGyVEwBY+fuSALzBJPvS/KhXt8ZeS1z
DTSEkAj+4OPZ0z4COH1oyNucvvXOayEqZrryLt07OlSUO0BBEeu0az6fyi4XXfU0QSdzvv0iWjYB
CxatG0Vqi9f0ut+leWKz1Ag8Iws/apXyjpRMllOe3bZjSCs00wUDCGUFj6JcVosj0LKp6JVq5PDC
bOxwszPZyZC4QUeiro1AM9bR7WRp0iD0gpoOu0eTuufceIG5EbxZQqRQhZsuBUXAtHJ7It2ae+H0
9nc5psSmqBp4pwHMmknzlBBkK7BBUXq2S4BDtqFP1EJZ5wjwogz0APCvtGFhwQvFeL8awq0cJBbf
pwEqWk3lvuWiXoHsLKiwkqTu7R0fCl16ZTcW6n/6WtMjr48Xyy2Z0j0Q96ltvZJeUYaQ0Hy8gK5p
Wiljfy/t6icezinvVm3PCvwm5RBx7sxdiOowjaxFrxWCBcn4V8zxHm7JEKWNiFBQAyfZeEAG6WSO
rtrVbuUliCqt/Slp5QJ+v5ds+iyPWQRUdvXLYQ22IV9IuI0fPu3bS4akuZlNWZyDhfH9YeUCllhT
A6PpUb7OI9ELkOHICfQt0JjGHT3lHix/ppJLNeXuJTwa31fBhkIt2kRwz//cRH+I7Hh0+7hVQHvx
gxHd5WiJGWVCX3Szwop+ePJxMCpCKyNzg8F4pXgoF+YftK+A5w6ZQsNvkq+t4rxGWBZvI3o8gf7y
dGO3lP8LXcOgRCqcTZusVv7tBtHjgWepMOoK1QQkdHwVNT+r5iTRkG6f0SXahA2tP07fcJwasb+i
yzACFv1ZvwFoWnOpsG0g08pQNJOYylD9Rs24JCWtFKNQtYWPKZn319Q24j8xMwztKGbwxfoiNzcv
g83er0EA/7LLyyhCRHIUnWpoY53hXbs0Su9xZURt6TcpoYsABHFWtMGu0c0IpkJnX9XDH50YTOPc
0kHdB/X62MSZTQC3QtJQwdKOYMaYrk8fCYtP3Miv2rfmlQziSVyMqKYUHw18PyysP8EdmzOKZoMG
8SOatEQr4/k/yfwd5CPexHqVv8bDm8gjZO/2cYolJYA0dd1/J4ppOSeAxZcXwZ51S4EjwoUaNtFK
EC3axSmil1fRWVUENWLsCNvEgOuh8/A+VSMbmp7307Fo9kbPEq2wRAO4CsrwOdBnlHusT5hfheXl
J/xSe7Yoj/hV7lJ4Na81ISBmjtTDeEYe2LsozLWO/eK9xu2BneVKoALvYjkNRSPzhxgq9G92QGaL
/ZmSHJuBUyV6mL40MCCz8BOkxjHKEuRJ4VEk7px0JHv6+pQIUWpzq2/dYaUAaRXr+xIxAIOeKujk
gLmOPIDvDxvbiiNMraGHx/L/smghNw6VoekGMTaCjtqmOP8d0n2oMPdbVjs8lxI6vGZS06QnRZf9
eyMRdogRqQERkW6AN6bDG0FSQVhAOFlf1iFTS+1QgSP3bUlKDa+uJFz4LasKSmoinNmKgHV9kl9b
IKNfTDWrmvThde4nsG8dufD28lI8sZMXknA+F0hwju4quZj/iIsVFoasYHwtXrjeoQMeUgsx/pAD
TvJciq6ZppIjoxqzqp3yRheZdG3kof1ztBCDUNRYcRlR1Elz4Keeat6GM60hVtWN3ibSFqqj2o//
3ouG2qZyOL3Rc4PHd+rqKWsuHjfyYWqOjo1XxgjzKqM4sqtSNlaLL38nFkfFDIOhZl6dTrJbHatw
47Gy2tSjaK27I9w1pPvx4y+vevSLCjigZX2Kvin1GOvGbtrteJrOVOyqCe3QuD+PU9cM+wh4MWJu
FsgM3QWrIDFqyy7462MwAr4nGRCvXoNhEKp2fkEpI5vqZ+f3nZq5hM1RxPiZQ+X7AhEhjkTuLFoZ
DrV1nlz20xAjw2j+4+BbhDt0ab9SIxJYxlwpi32ayNnAJ5xj11i1KdybsjZ1SBq8J9GMqyotjHms
+qrVZ94Vdk1sAF/cPphibr3BMOCVAlVNwc5ny2woAQMeA9vzXsKdKg2cj3LecYdsoalbIveY4rMV
Q1gz2Km8heNhJJUlTmJSXhQzYT1YUqfWwJS1qCYlt/edfhwMGe75oM4nqZq5yH/arMRSmfpDoMYv
NvopPzLyKxROoDZgV8amFo0MJumcPpqKE5hfKQnCbUZavo96Lc4ynvZqPAdedj7f5scb6YqoGkr3
2kUx8PeOkHOxccGvjEcHxOzW6SSNuBkY+B+qPFsZtcCMtDrgCGm3YX38u9s8w11pZ7t1Q5LZTcNw
7rHgcn109zcuk3KnChbFhiJ39hK7xFlFKvlc4ourN5Rv4MZOiFnO8/frJo1K05KzHrF/QQhR680q
HbyudIqN+g2wlUPDBDZBQEpRUPWiGH9ovSf7givVxQaJegdwvXmuArGS4ylJ/48Xh/Pen/vNL6ce
qksUcXEgNZ7I63lhFcTOB/8ftxWw9pXVK9pDefZNt6NVEr5ZbrdPovIQwRbP3D0VRud589WlClTA
91WlLTZN1b6horWIBLinjpiB7XelcukvBHkN8xrDIqgcP/5sCnu179wN8ZmawDFevsFrbg+sGYI8
MkH5HDHzwufByok1U+II5KtiUB3iZA2QlDYjB5IbhyZOgskvDPo9y5yeWQYej+YcPR8/YjunnDYy
t+GnHhGgkRkEQmPvzp/B1izVIIMCXuCIa/nJWFf3X855hd7Iwb/Rstru/E9BKnOeKsC0a1Zxs9ut
Uq3e8jJ9mDOYNObvjLeiYEnua47pxCtN1dGcdwtzjy8xB6MPCFi5WYlz3k+8fWnvLBEHbwsHuK7g
BiR0/CYprY0qfNSQY/CEJJMBi64NApTBesTKWhRK02JT5YfKoMolrNwsDy7SvV2ZjGZdXKN37owx
jH3ikv1GIAXGx23pxSIx9ikh8ovTy7LQfvyzFz+U9nvlUOiYn68chOuSnVXH828ceKw7q4QWcN8T
sUBe1mHyD/xtx8cAKW7bQGxj1/KdK0e4XxVBHEWmRH36UyYEYXPHv5bJC6zKMOd6NEBcqmOklh6Y
pvD4XSONg0AxlTORH7NVAp+FvQZDer/5TZE7h16+Es3dJqnDLMxua7NeImvQbHaKkP3Z+0ukKy1W
34DcIIJtXuc8cCHkVk2QLl0bjgb5PWsw71KKXIxiitxJe6CMs4NDwLASVN4/c8XVK27OQF+C1NWN
pp3z9GqJtTStT76QzfNq5G3fuHdRnUf6UrD++81XdSCBW1mJINwhYslWtJsltgFr2MY8xzw147kI
Kz4KKl2L1VRHezfLPSlnzykAnmHf9lCGAM7z+cy//sW/wbQ9mkCtRDZuyuNlfNMqBhoi2GhfXwVD
UCOHrvh9AD98K0FLSG7hUEKPoQm6X0Jup4pjWv+jPnAzKXeuSAyEUTrurIwvgt0FeOFsOdP77Zo1
BxXs7iQGzwXE6sl5/zQs48v/murHevWQBgLpR7d81hS1jhqYTJuA3FpMqx5C051XGBuMOnL6HIw9
IybJYHaCqDHTOdopo2TZTITwwoi85EeMzaA2OoaX8J7UvVpkMKlTbSfD24vunATnb+ro8zHNfIkK
nBr1Zt4XvOYsVltIdw+OIajEop9AMeANHaTsqSamWLjoBgJP9aavZXIL4cKvaXnVXTmVB+cOsp9b
pfSOkIhrj+5DiHvHAB0j+yfx4Xg/+qwuX74cjHSJZzqLdDhAjqAk9E3gLD+/f0ZunMssvu4Fe9j9
6MZ3DT3mclojE8PocwFV6ZprsxlUesk+Nt5mBFon6fEiNYchIR8mipPFGgE7zvTOALA0vpVhN/+i
qcfaLJkCQLxW1aqWQXPqV1iNiOEEbEOtBEiyHDvXkW2ZHjsLXQJ7Qdruqu5UAUCBjGGRC+rj01DX
77yKGxi9gKzVCoeVHdSfyXE7aqyJtKlE1mFPpDP/wd8Bs/qi2KnMPMXH7sOGTObp8kOX6+A/8lX5
W+olf2vo/3XbtlL9K7D0vbeSmi6PwKPCByVaWWppAGEihjyMqnPBEAM0WLowezOGqS08G2SqzCuN
YMYZ1yDL3t9nYjkEwjIUIlXu3X8sJ3PU/0SDvc8IO60VickHUjnrC79LzLxxleTOTWZ5beHHZ+8y
teKJzLKLq17kCWzmjqZ9JmuFnzIzKXKSX6X2iusevvEJrBV+FGDXjskWMezA+kpCQeFKFFfvLEvG
WJEHyH2fpnXmYDvyysnpf89sMzeTIOYQFRs0JYhkxYe7jbvK/ecNfu5twebuqZq3/CaO0UWM5OG4
E0qXncS5js9eHBQk0xwc0gIDg/T75VvoR4Kl2zimUEuej8B58964ospdtXDqCSJyyK3pyoegjj0e
ArMmmJjmOx5L5jIrzXF2QfKm1OzWeo2CJoaqdvR69PTMzsUbyePKCSgQu4mLGUxH/z3SR8majRKc
QgwWmsQcoo1Tm0TR2K5XDi9rjpHDVsKGAjH6In33lgUBKOFiX5oo3iN/eWBUcjRq32SKPyTyTxVB
PYnKB2O/m/YbXKcCl7qlBYGZjSCpVIbjxOOogvybooNx27XnJkJvnli//hyDCMvbM14RVrT5lB0j
7NdSyZSCkOxYu6wzrj3zfdNwxtXLMJ5LTilpAO8G0ia88iJNM5LM8UUCDfWEvr1j6283wZIURd5a
ZJrd4ICbUts2pe4FTpUdCOE/DqJZ8EllLxmkSDr+x7gJD7pagvpIrisvL0XK86YukY5IH4HqZGyS
AEvsFeOCls/mNqUcVpEGElpbZdjPcs8JdfaMHSBCgzUb4HG1hjwhSTtFAYEa2BPYJPyCVUzioA+A
OtgvXFuBGO6SexOKwClBJuF+v5mpaQw/R442MHOoL0XUzSBDVoqz1x3wB2itgkFM95HityNUJi+4
/j2gAr00NJZX9GKLYigYVge8I/QAPDysBg1/jzZ29rnzxpwmAvBlEnYUHZ/lhQp9khkNM83CKgTy
IhU6rSeYhwNw/IttN1569m6muLlOi3ivIqF7lr8ubfXbTWG+Rk7LnBnGN7XEjj0k7lycEAYCq/PE
noGlmsPPwEgtJIY0ciPNcfaDs91Bitb57RpeszvjQU3Mm9pBcPfrbLbhjAfLL0B6HVELgExnOQCS
VMEhIUUpzEGvP65UOGsNGmWvVdo+VgS2FIbAttBazGhXfdyiC978wtI/8nxZDrfIQn3VLKVJs0J3
pdKlO+nX5vPXvP6uf7KiyueRU5gfg0xYPjSGqcEgO8QUd/WIldJj3THXsYb6/V0mzSaHGxuurNZj
gbmQldqIfkn16Hc3AL0TiyuUrMaETNndWLNtkx+iNSIXTOHt1L3QbcXFcBuvPqn0/iLSOb6sCrrz
QhK+6YRFIk0tdfz5gDsc98PF9WD+kkcOp0svskcChKHK33lGrwl+rSihqPxGT6GQGPna8GXomLUO
z7ZSpxmDNsAzECLJp8j5VT2vzB4901Nd4QDcCjhrUkCPNszYqUccwdq3Bz2jmgKvnik3If8jMJyJ
aL5yYGn69A+QFMyeN0AjaL761lht21LS5/YVIMtHAy9raJeF0kxRGWvCxdY0iqHvEVdG3w6lw1v+
PolvNLFrmWaa1HdLdekUGvZHGPU5Sb4dN6t4jBBbTiQuw7dvni9LM09dGYWiGM4JPQc4EhDbTa75
i4pC95i4EisQnhK6hDNFLuzM+5+pZZF6KQnztLdA3VjIQuPrH3hpJloNmoQ8+EzpjhTxDO1JGH1U
Mj1mRHbxa38o/KPv64UaOsp3M0xsXQZ9nN8Z8m8gmQdjUeWF9JG5hdq9q2GyNye/NLcE42C9VzA6
C4cHem0V5B6vo8ubHYDCOUbLwmLfzzyfOSBbxrHDSuzZ5drSH/Z56/4wrssDXG46LexmgihQex9b
Zm4rntpvgN4g9ZHbjt32a06CY/F7WDKGm2+wySnnu5ROZS5hzyYyvpZsj0toKDsUibrTzdkQQwd3
EGVIfJIeXq0vGhQNfEbJIav0VEEc0D9YThzzcn56FlAztX+j4QsdC1e9ZGFL/P0sQlR+UlWxm5WC
WAbbwOXEkD/+cNHXAy5wyYEEUhaUmG2/DD39W3GToo8fGl16B/zodNEi5K7iBU5URt9xwUp/3Gf1
S/I3cHWrPHG0yKgg+V367gDsAkXps3iY4gp2HS1V9KWO9ASzmI9boyglDNlhmbIpGfWDRx9gnC1O
D71CiqJ83FVi9rmfGIrdvzW5QMEYtGKrYT7C5odsMO5/pFHD6+zflDFwoBFGBwZn6VcsLHufbxFp
tJdH3AqSOe/qotrgRq/Bb2bBQQRj0vGuxwy79WWE3zm9JCMfxzihNXdyxogusht169QYLcL9n6Zx
+MZxng8tLOYBeoFU4tEBpyqWKUIS+Gr/G5rM2J5ZbqEXNrvD+mvl7w1gylo30WhP9N8Eeeqmx9dV
u+0CWcaX8pMdB1RS6o9F8SBmHVOgqgJqBb3+mbxH8J6Gr8K4plcTZ7hDVLNj8Du3XcivSi8RdR0s
+Tr8GNXTFVEx2UWP7fsq1F5CxfuH/qbaYGLCPJvd2gGkayQNfQUCV+dox7BJBCw9yefAQG7Td3zu
uTvR0giHXIqCFvFPtEvdXFUu29uOPDYxDcUiu0KRADa/YbQtZzLTYshEoPpO4d7Kf5ilDvqL3rDk
hMY7XN+C4RFjdvD/67qg8Ojc0guGHF+JVx5RqrGv5b5RHZQrTiNyA+KovGkhwtdO6xRYxArMkCnO
qzb+UfALUPEyO+opN1ktHVCnOtR8vSbR+xxzXqRfEWjztw09FSSqlwxlplLhyDYUvCxvIZMZHTv8
NSRt1XQKMu+1gjXs/KzC/hOrQGZTVB8pAbn7yHvCYOdeO3YwCa02KXDdYp1wWE9u5K9Xgn5vX9rC
ZAtZNitpU9i7ShoRvEoeN5FhaMtGjLxcWhm/lEBe36kft32vzG1T/Whs05tjI805tXdC/q/AKE9A
ipQ760+pxSGl2MGVuTtvjxFvwmBucTZoN3FRDHc64nPfdtjVpBS65wPu0Zz+ukyia9RL6YhTMSDm
8Ylxk/m9udiQu38LGvld/9SF/RtBsXv/9tPezdX5FliE2voX7j6sXG1GRWeFNwTSFbrTt08huMN2
29GugC+J2qKQC9WH4s/0kBOaPLXNiMRRt1p7/NQYcH8hIJvzeSq0Nmk4fZXc02lGmOUfd1fT9/1A
1CSxVuzPnYGOjpWFEpRBVEy5yImxHhwztNlfStNsSbeUaLGCCgphJ3xRu4T6RFHl63hQhVSUmQga
414ORYOMo5y214ISTW+b4wFk2ciLHPSBsrE3citPx07yBhfG1Z02FlznDWjulTCFB8OuYmCx+xBa
+YjZuBQ0eMXilR3FvG2+Q03oPq8kHidh6YnDDrxI+RpremHToKrMpt9mGyleoknTM6r7Bq7fA8Tb
qJ3HA+liTfXXx4AwrXw+N8ndhzCw+sGCtZd0kSq6BN8T3QlVqG2bpaaNQcq+3GN2sGPVBOZC6zmZ
AO9pVAV3shFjnLRym414NnrhtAl0SwvVcShDa76PTm+jRzjJoPe/r2cwPsh+K3O9/XWTuSH2HfXM
1Ejpdur7iCfZt05cEPR+rMcVKHLYB1jZvjLb0uJCV6s+I+pvTOTz2Vqq4cjy6LdykoTsQOb6z0X3
9fQXDiR0IjMPkt0GlK53G2v3ZYiBzSF1Q+WxYKIVS5oH9AOWx66WGy9SqIN/nmwZt9zJr3zB4Duy
QMtHQr1rxZbEQNr+0Ziffy+LtAATgXhr2G4cME9nReT1/e9tQ7bF7R4+rnZ2qGIT47fgIMHdDzEk
uLqZhdiUmnYho2qvRdonFFqfVFgWb96OJGgt4RgZwdbmoc35S+bU6WLemrYHqMavnTxDWbp+IHl+
6B5w4OsdYmEapNvPx+zPDFJoMvbcbOcpco999tOsTHtGvNkSvAxnO8w7DVfeRP/IhR6hGvVLy2OY
A1ZVb7lXpCRI2ETPoxpIyIeqMaDzcnrgieeXl1JHYGFf1yCXWMjxi4E1GEL0/2Ngy1CW/++cVIwM
nvJkoE0b5mtNnFJJhtcV2Ntvm6hagCVTbyM6AMppXTSajlwI+ZQEOoz4SMN+FYXgti4zBafm4Uw0
7fd96Lgm2SR+EaQ0wFqRmaWdPUnPSMjVlK08tv8sqOF7ini40mzSQSsU3+gTFoFt59RaCWZvlvZk
Y70z0aZaUnW6V6faphkKrOaI3fO7bzZTEydyJHVpuidVxhcjpMa7G3KxRhRGKz3DowxEb+1dvDG2
N6uSPpKjmamomsBTOqFLR9lF/gzvjRkYBmKuBuqvnGGh3+iRtwiUylbnAJJge7mjXCY8aqMeG2OY
5utNawzapdVOIUBD9FWiQ6pnpbo/+zep2kxeNwR7bRjSdjRG4/6eWjG1psj60HVq9d8+EzHHpdDu
AIvcmT6y4psvXdgCRKolGp3ZDFwDa1/idxUSQcj0bjNShAoVWv2oZzEttVk1wUCHxYHyCXYOVNz4
FiFW4dNbPA0/A1e+ni8RF58Gu7CPuFkglAMaSzbbOmawPCXXd5cOHJd5yaM/HFZHeO5L075EJXCp
9lKfSkMfqy7cECRQOAiJUQst50xhqaV5bhYL/FN20CCQTRSMytM+v8PZt2I/ACR+eWrB0cQjc/mR
KKbHAtyHa2WRstfySR4+lH9FWI5yXR/wCcoxMgcwwv11V1TSw0XD/aN8DIKD3dJteCreyZPAz3GN
UebGtv18vupA416ZW8kO21dfvHV78WtkVZzgohhOg6wPjkjlmohqEPEdaVrPZdLUWZdYUTgtPm8D
3B4CPB6RwrkBZFysh4h+rgEGTAlAPxQZX6bwZCb5yC/DVAM8zMgHYVE3W04Ui39iFxycdYvvVb19
8LGblFIL8rOCDiKEvoc85BDYvXPQvRjssOQvqh20O0ltivkPWrjTNUMojtsk8WL749/OOSJAFVj4
Zl9E1GC+qfRE3R5Zm2vttp7qxqamCEBMiEIQ1oRSvdnWDuiQIilLG2Sz3cGSvhXjMsN+hbrTRnQj
bW98pZJtX0Inz1hxuksylbOACImEyfCMz1hac4VhLr42B49xCJ0PD1i42OAwtamQaoWLjO8qcgmB
1sD7Y1Zbw928c/vMHGkQPtuix5SodxO1YYuktMDdvdO2P2islQmLDKUvZ5/uxFuv4i0g0VfPaEXN
Ihxf27iHv2/fLbhxb+aH++0um1ZluuSDQ1vuzjneifuLSVGvipl1OVSQdJfqFmfGf7mCsgnakKYs
RccQQee5+1eV6FVp+tSSUVRHbGvphJZrWhAgk6Q3n3BcDxcZkRpRlkIY+TOqScCZ7GM6ztM9GdPY
tvH0hj4A3cZUOrEsC0zwJVHp1SweBv1Gfo6DIERlZInY8VkIqRVtCdkucCrGNuluN7rWvQnMo89k
N1DlNA0VN6FMBoiqlLiMsyUM0BCbiBlIgEAByHv/JjT4sh0BvkP3bBVh9G5YxdymPlV1VSHKeKu0
KSxJ8mrml80F08IXEqMSA+llyNES4ES9CvBb0YQf8gDvv+fsgSCMmyBal4RccGtlXy7XeOW2Dmas
Ir80dc592RIsWjJXrI6FaylMp6Lac7/B68DiVWU68llx+WQrKsXntd5vkRnTBELFNYZ3KKuxff2h
C3ye2GGtVAXYHkUBxtX0r0rAtl6BkwJik/TAcuksiKq4u12NmYnkbTU5KHBKer+EmLLCv5JRR5Ob
4v03HYpXlM0S9eGIRr0B0t0SwW8if4V3KnXa3l9pYxQ4fRgQOfwSN6D8f36cZZsGF3WCnh9X6d6T
c7dyRM/pVnXyl2kwojPbmZelAWPKKCEkapAqWUgt/0EfjBc0GOzb8lVtDcUkZ86xmQbZ85BibcZe
SFtOeFWZ55kWC/g5FQA5xIgd0NQRLsVOODwB8rIdAZR4PDvLnE1BFdZ2AQ/Qmgfj6xTGdpBHHWm1
eA8rsIASKd0qBBtawL/4I0pBzy4uMQNql6ntORVEQ7yU0jS8eYD9AIdvrEQtIhTUK7uW84+Jz8zq
qyK7a4hFqAxa1pkowQv6ZkwJDhGam6eRGp4J5UVdZ+Si2WuZ4iQMvQXs9iK57RJKmw7T26Xqf/Uq
sQLZza8tijTsu2mMH/znPbTAqykLLdB8eVtN6No+NNDEH7Sh0fay2hs1xTXzEWK9HLeuAoM7ZoWJ
lbsZjNVmL4+ykr9lt2Uw1fEAnrT9ypww55hH7+FNmASLpQOS6sRvgUoTPPyb8G3IvQwbshcD6V5o
vsMk4PVM11INW8eZj1k6A/WIOy5F90o6ZL/eBajqM+R0V0miFcVKx1PXnQWAR7a1zVYJ7OSuMBYl
3/tbu+lvkPg+PO8dzc5fYlTg4bggJkE9xDsrOKNNcVcgwN4ZCdP+F3X/ihPy1pkay/4PgdQtrXK/
LNj2r47dnLVMAq44RMcUC3GhjAxWpnaKscxUMkimIpYmqYEl87WwjYZxRCzC76KhGZNqI+cIBfBz
9pEapV+9tHD6LQ9FITWwNfWSQvAQRu6Ii0F5Tsb9B7OQHZAaTOOGvcAkKyIWVS6ltkYpKGiIF4h/
4C429IMOv2hN5o8D5jZcG5N+PMIjYY6NvGjr62QOS42EKbkdMLLYAQtJtb8L+hDG8hTSnmz+1cKt
CNPWuhvA6RDv8rvy6pALKs9d3/Ljpvr9j9GDpn0TuFWOkLl8bnEL+yUo5qzeQHMCxMHrn3myPkuf
dcNAnxqbc8LgSe7/EmolAVYzIg1SJ3S0SZ9ctJdbvL2a2ktQ/2lNmyRo6uqlZX1zF+g5KcZmw3lS
GHWfof4fB2jHO8oxxLYxbt50G/QgKqlUB+nQHQ4hdrCBZrkwR8OxiMojL0d74KeABJvqoXUzxE+Z
fRvZPjAH1pWTMNaxOoAmVzRpoJ2k5KIQsqWPwMhrs52bQ7AAODvoXjmYc2kgZR5w6z8Gpk8kJPei
ZlIPcN6zvnwOsyto5OJATS6Kg/emQqykT69Yo2mzNB0/2HO9hbWh5i8gI49vn84UVzo9a+DQexnO
ElRtt4JoWfUg6CybWpR2lC5n4RdPjba7uy9ezY1/jdVRB2W2U0z5T+87DrO0sglvNU9E6fotcjR0
fcbUxqUI3IeBNeLWjVokioJ89gPdORL8cgOLrmyzewoseXqVIWLB1Vck6gmNp0rpd3KFrGnSI7aa
xbv0pKaSwDVPpsdByXraXEUTDeSdoabuVK3HNT7L/mrt7KtN5lo07gtr4mFrkB5t7dc/je8pfBme
BjFCceTxCGCLJvAZJHExxMojMSz7ZYiW3MWwhnH4CviHUKZO2sKvSd8YlLFks9OIOs/yK3lWaHCL
+eCO31e5QAkZoiVmT/R+hU8W5KLxlYYRrg2OkjenLgr2QFEHKpx6BBAxdmuYFo87f5JbG6INIL6Y
liqvfbR/Ge39SYp+J7aPvP2vi0B1jJXU2aZg74rw9ZRCbxx85dQttFWauAChOwOCYColXH2AOFFD
eEHeXoZs8PreZHvyjVy0q1TZ6cLUp+uCYeg8rC0K2d478nSjDmyvR5xnhaoWLvXGYxkr4tpePV5s
M/KH2gboMJ3GcnsUe1rkyYxEhiHZ/UjKcZ7Bc3ujI2bxuG/G2p9YQtOdusj+ZKoFwZEQwFYjtc5Y
7iuq8GwqztSnu8CZRv7ujYkLphOcDjTt2ZHTgAQl5C7Wx0gMFYXPDiWCodDdYvXmMx2KTXqEormB
+XN9c+VN8FjQj5m63gDivmMnH1qpKsJoMbv9iQbATXt41KpppOEyEFDKtIe1MpaNTmue8FLVG0Gs
kRORmdrJQlv+gY79ZC9NUm2zH73HO+LbZ0An2CngEXoUWuDFM2bKlYxsYbbGNPLAliQz83Lrqw0s
plGq2UEMrRMMnMZbbBGF20vCwZw1pEnBXGLHyp9qn5YvdR1rtF8bdDYt+IRGxw//f+Y50wrmGA5i
5joKWEGsEaEjdH+p7c3bMSPe81cFMiVxyamfFEwlUGSEzuqQXNMmK0/dUqs1ngujjIedYMFV52Xh
4LS+oq/SLD4KhUxMMfesN3IOHm1VjZc5/DTFzhVxuHbGRjDsbzasdxh+jX/To/k+HsqL9arhpql7
bvCqog9AmXtyU7TXPRbp5m9Qnw3quNzZHHf56WxNXtBQ1CnVhGx97jxaTGQ5MyBK6MjZUXsAjn8A
zLXjeXnwdEpWiACPIfvBIZNgNTGX3h55GpLCSunQq8H3XDCraWaqVYUZ3Pz/Nod8147dVPlXGuQF
qTxrNs3ez+RBe2Jgk93+yZ6hdkbvgxg5GMPh+d8aF3gUpIdAkZ/4wJEoXsaa4vXPQt6ZijkESjRV
kKkq7mjg0EJGVSOaUKD2baz/Ejmu2mxS+9A3/X3zGx7AH8dvQgRsqDRYanEN8XSd+ZZEzv5mhCj8
HLC4LVoDlE/6+ySFm/z5xkrPfe54kZefESqzAcBnFNnb2rmGE1T4y0qEhGcz58PpQqi64sbkK6XZ
VVdLZ3gqeNcK8DhItwY0WpCnrewI+45HFJjRLWHc5TLMAGiL/WS5P9OF3ZtsB7HjyY0m/tFK+KKb
BiTtJQelaaK5L9iGv1pI7JZfOMsdAEcVpMHxKFtiF5aNBLBoij2EeZRNIbt0Vy1qRuMxXWnRf54S
BQfHp+SXn06LnY2ZVNBFbbkB+t6fkVKla9/qx1qbKVwGgN3tLGALU9W734IppPzPIPmBEtF0/Zgh
RW+2OwycEHvJwu65zGRWu9NzQx7AlPdwzGwl0U2w7u4s7hWzSJZeHAX70mjww5qYNCX1NMh00Qyu
6r/o/t/m0uDseDuBy0k0pQeKq24al0E/H5eT8fRFECGDaCwO9QjwuS3aQltk0KwitrZFmyyp28Bq
5S7Hd3BtP4hgylH+1KE6ZnkmheaixOersTjHXukf9ZqDw+FVv9muKtTgX26mibiR1mT9QuSgEtub
A/7KquXoCbxQb138Tkpz/4k0cyF7IIezJ7L4e5weyIk+LzO7W4J6fFw3MWy1IKBDnw7gqO9T0AzS
pbMu2g0wOZbN/pQ0pnBz4SsbsgXaf4Ml0toWTE22ByfB0h01TtNyJyA7pAt88XnXMI7q8CnPLSRq
zjhJfuR8btTd2mB+3EOT5xNO0jjFCt8IlgliU/FeXKZMni7vbTo8zhl73tTXlsbshM42al0qZq+5
pBYcgCnNTSa8p7ZgPJd2OZ8K0yCm6PnUxyBEJn/K1wWgiqHDDvUxbaU/lLerJREnzcFtRAsnqc25
CwbH5Q3dmdVS+mRxhWVqhHL/l1RNpCQEhMPkVsa87pLk1OlJzCStr6pLUlZv2ETguXjDhNRGyphF
SaYhlSu8ZI6FuZrcEVEqkPpNHaOdanpQVYLDIhdo342JdMorR75Bb0fmYG21OWH1s3en7wLeuGuY
MMDg1/7120J4UJeMey5g5xA0RoYyEFMNogrBHp6Ot8+T1+gtM6IL8zKKhOhEpqFwdHuOH3nszdqH
rJm6BHKHp5RigHq3j5quM2qFIvnk2357tTp+XuPiimP8Md5fd3dtUNahW+GizZtM2l8Qq0H/55OL
kZxzvkl1p9hYsDCB0tUhRiCKzYRA0VM837RJHsyig+fMwPgEp1YknWg/ST0Cwkye6VF7I85M+B7m
2qctaVnNFjRLOj+lcKoYYIjPmIVgBCIbKV0fnOo6qQP5Mf2PA3fYd7p8LCRJDHZLRJbdVStFvg06
0WKnK/ZmKHAj8st4sIjT3HcNFenT4PG2eHkrRaSmWa/sOB3LmMFp19f4/fy7rBek84vkKhqIuCH9
T68fkql5XqlAuLkjUKycnZslIuIB6Mbw+MdEmu9Mwt1zj7/+GF7yxximpzqPm4LaG02UTDP0l3rd
xdL/+U08rB6U2CiOI6PE2cZQ1oBmaKAAmnI9SS4FxiQGHL1FaD9KlP7BZk4Ar7CQ/by97f0cdvYy
8hgH5/bJ0/jyleB3aLlmigaBOWOmcEMprecudyXUMH3Fr5XLZBVhdT5JCk3Ssvk6TmwVLnq1Rkfq
dD4RRUeveuxcX2Nw1d0CWD+p6dLlUJzQPIvSOBUFmwYrbWMrhjT3XCsjB47XOVmtraEE6ssBcohn
ij22NrrfMF5E2FGdylHVCKYrsdhMfcQ9lSCTxr4nRbGecUi6Xid2HJRhnh07w2+d80GTLaCodhTU
rs4Ly7B52FzVyCu+dsoFKVyjjEohYGXEduPaj1tzHabkQK8sXVWTnRasbKuwrFdmcLcJtkdoXbdy
+e2HsKQRRLASrgaiORq+WCkyzQu7ac5IdP1C5WsR+RhaZoXpF/qm35W8xPo11WZ1j3Y5qicxNjmb
ZJYPGNJbR/lpdZejQCrzZ0RISOG2UxdULRP3fsTgwSTEA+b84DdIEzW1X6WUIfeCjdLuwuatorqP
rc0DGiFDnx1aCumkp0f0OgTCXZwZ2dyH2ZwgvWkvR9SEFU8MnNiBQO3/goaMvUzAOOq2h/33ONWY
80RDLsxdWYtX91ckPy1/iiXAUR84yqHWlji/lHiQN4a/9+noJEruEzdhSHhew3QzzRG+bcuxm5tR
YduYyUATsI5dv2iJQ5BLu4RDjyzyY8OVxOxLWAYT6EGI7SSeH6A0LfTfPQqx9kktSKXKoDWzAJuk
wN1fNdOQSJITv7wXlCCQHBjZrrHuxxaVEjBcO9jAByqRMy34qEnty0wxo57BXDbxKDJclukZQi8e
WtTSugZ0xwtbkzld5WCWcBAApBKznftkRbB+1WJAjrKT2WTAhN1OFddgKckQHIGwJcEOUhSjxL2M
4g90ACHLtgYgftsNoTn+PvrwaXlEilpmSO20VQQteyS2VafmmfWOstaJMweNyI3iSnzsWhTilYJA
PaWlXDVj9XhL/lEbkvLlvYoPqjuDeFNVQsQsBOWITw4U4S7xjvEw8Qp782u46oA7DVsjEN4YYAJZ
Vb8qkS0SJ3AM+w6CqBCv5hFPhypYrpmXtzOJ9oqnxmk+8ZqTQdHj16pO2/lDFIXinnlmSUNfjFVO
8rGbbPQv0IE855qIdM/5QzCCBSlSG+ro1Z/ZcDRZqRpHiXw8i5O1hxiuJ907DDXHhOY7FXgqgF4l
cu1TazXc0WQc+I4P348bjmvtkADrEPXbsOx3GbdvJ0nYPvUziq0xzC+3AamOJbatZbCQ1XT9WEu/
dQ0QGR2okF4K4GRJd0rcYvX6oINitAWy1LsY09uR01RUoVFNtPcL+A97meDWMAPRykRzPc5HGyct
aC3YxK+KC7ByQGImUs+RqikanONeGOsD1TPfydgehdm6ozHO5LupygQKdVWU/BGbVndaNBNzuykt
APFtmgJnSIrpn46GOODKU5rrHQkPZqy3GyDO7qlAMeyrSw464ttAe3GolswqYkj4NQnwZiqvmcgI
JaDhp88vDpLjiaJHnFqXqLyA302aVTvXa9IoisnlEnDp3ylP6Y6n6mRNwUXh5NSrN3J2ijjYgCic
LW/t0eBSS4DLgQRkJ6pfq2lEBsQjiJu87mDNk3E7KZCmhk+O5xaxtZUxDYNgcEYEQ2ogY4fCoZPM
b2edyFC2/f8P4vMUwXlHulhvKoGQeSguANOhohtPUgMlMemvCBGF1L1/TojyfQznLZDphNv2pcQk
ud1b1uMC00NqCIKeNyF8qy5HL+Eax3K4hgxynB2a3v4Q0odTaeAEDnVKXuyf5VFUKiUrTn11S/K4
5iqaiEcxIlDYsVdZNMEDK7QTDdqich5pMnnMmXeQ+TjjBo8Xe5NzjneEYo+KrvMb6gFY+eT+USj/
35PQ+68iCYpz/QdKnoD/rTjc+2Bb7OKKgq0k1LmQC7rD3MwRRMsL/ieoEc6uT5HUX67Jw7M6dbQ+
nhx+nYOapN3yFrLrvT+iELv6A+ssVtANNgVk5lJBBke5nTloKKZKUqtrpDE7MD8NCYna8kQpiRhk
mhSDDWONZin5RA0gL8zlu5Z6IJ/VHGB4CrNBImAIMS9+5adgSLKwYg9CFxf9NFjV6bfOjIzPULBh
RysqZrnIHBLNGWczP+NqfYHR2jvPhJmC6ioFsromj7W+J/4KmNXFXnt7RqTN5TKEAtX/Lxqt9fXf
qtwLtkd9ubnOwe4Lx617dqSmSGeIQ93Ej+ku4Fncwc4WsTs2i0B6jDj96ddiiPqreDa7WA4HaFzq
O52MQohTtHP7ZL0IMotn7nsmkfS/qvGH+RXo9QdJf1AHj25nkT0bwVpcLmRdGJp79MjpFZnixcxy
qNw8mFqlOYi2DM2Re2BfYphJCMjEW1zBU0kKmbh5XPj44Kbh6noyg3G3Oa/GxDHUPhnIJWa7bp1x
VCUCwSlZPXfy08DuIlAeN6rFzPzVlVyIJnmOdyBXZcY2Jlj0JRTTK7GtUNBunU83RNfGKMqnU/x9
u24YgmwwxoRXliw34sV/jzzNFyWZ+fhdIdblOAsDntXZw4AzLQL0pkc6RJaQ9rbetPCt4HctdSKl
DccWV/YAjeJp3ofDb7Pd5bp9ar5yxsJpIDUbXGG2ke214ZyEOlGN1sAJiC4x4MnZm9PxA8EgKSt2
H2i+R/rEICIL1BsG8HNdHgfJhzaBKP3gjSFvZ8SUMgrTU7PUJUa911rQ6JPiNC4fIhOB3WyhN/Jb
XUhX/6BEH4cAQL8D0ol6tznPNJlzqbNTzZb2CRt63srmWNvlAZztSOE6bvjd/j1D2+hdQ9PgcY+q
WjMqUrMdFWrLu/TeszE+hVEqcoHzWBwrP4vVeHW16EpYJh7UfRtJBK94LZtpRAZ2WKsBluI/AJeM
L1g+Bn36O0Dw7+bAZOkwgFKjt4gmENzO8PnuWURYpkw8BowzhwT2XFTFUTZJqs7GsrsLSzFhShKn
1Se53KvY30889ZcCDfHkOyqv0hEwgX6Mb+JiFaHFjMTqQyc2Ez/jmc1MN8gMOnZDF73afy/PIIoh
ZvP02YCVbZb1wcEBzHFlSJpifnwFmvlxDVGCdfchxKoRVgCtCA2FxUtlFoo01NLO0j0bIqBxDJqx
CSOxfEKuwFw2EZHGKr7SK52hyaxGJZkdaPOlxhGqdaIvPmXBlCIAsBn5HqLDGKmkoV3DixHgvylV
6rgLgTRgobpqRbLsjZSicC/Nmt3hYTkJskmYzsfUEIGtN7XWFtj5QoynqBrI5NOcUvJDJn/2aHFT
f2cigCpCVN3IZNUaoYxXbtnSVvOdMf0+b8nPNXsCTNjHiJvU/FOsdBKlFRx3G2p77DTXtIvFMaom
G4yXIz7utCitpSI1fOcrWTH9erVmgPV12dJmdR5JE9/o0Qw3hE7D8leK5o0Y9Ryh5ul+JCtHochL
hUtcZnsJjsVJ1RlQ/djr54EwtrfX0kdZGQuMHrIR6/dpAr4dBpmMQEv74HY19LbfFj3r/WfD5y3a
RZ9uPwVbvBocIaBcbPXLdva35+QZx9tem6gBMiFXfMmYh1h5Th5e3wk+l+XI2CjQhNlSGJtkiiuV
oArAduwjXty0hmK6GxmPPyhZ+uG0mWHmi+90Su2BCCDI6RAesJGgxHDlVsp4ewglKwmx0sS7Oqs9
236siH4BGHWBRMko7uVMjl3IVGg7kpZiR4FS8mFjjlMOS9NQIAobwX3apjSEL64ctQs2vJvAXeG0
Dm7KyPhLOtrvmnLKcL03UXpzWSOaxunQRiAsDcQgf5EPVkhPLXWn/m6z8xHIJMKyeYrUaa2XVJCX
CTqc/tH48iwslMHi2bAwJVHteTA2CUiGx8dV0WdFDJU9lUbu0U17HaeszDUzaMBoE2dkCZmXPJ7J
7CgFiLRj+IHac8WsAplOOofvwM6J61XRjR3RT0XJlMr9IdfMEeRUKMfuUO2pyozw06CQebjI/UAd
qv2bOqs/3FqlR8xt0FEijywHeMN4Ncr815HUjbme0CcA9u2CzZ6SPQ1hGwtGuCYhSUuW5W25Y33L
GDQj/TFbS8e1tj1l5J2Fn9hkRX9u63XA1VL338sYSuPV873qk/JpnDV1m0lxde1Nj+nUDkrYyn44
8phKc6rOzDyd3/DoooSfEy7N5TnHlxJ+3MRYkYEjWJ0VbJ0Ql2kKjdVEC75gUQf0lptBxxTR8cgs
JalBQor0FF6zNNj4WGvYOt0feK7Y8WmD2THZ5Wvt68L8HTdNiGzgFpj88NCxHXkt5GvAU3Gt/9MQ
c6O9ITwsU9FOOE8FmNREef5LX7CEp4Dj2n9qmVCAAWjmgaxTLAX5jvZ6lYASvgZGgXaT4P3KfJMy
NOIef+Dk/ycPWyqN3BqEUmO8hnyzeblwaKBNLilmENj9iqrp2DfBpHxJ7HH8heuh2r2LVcgzrbfT
ZHQtOe4v2+FIukr2vj4/QbGkncrrExantY3kH++Dc4WXhf8qKsN2y4nPNHREIdTIaLMEFhCOQecF
ALeBExMAzmIJk3MRNU0uQl3liccZ1QkwVnnG6shhAGQzGOsFY2eOe3Rj0zfFfOylBcIltiLSanlz
QyQ1Ycb3wdyPebbnw7rGhDlnp6wY4ZSxrcNo1u6mKqssbEAWxSfF/mCx7ZMzPh/wkJbYRMjhfwJv
DmMwjZvI0gETA4FZIO9Hb7w9uJlKZTfaAVNU+3xn6GT6PBuzVyhT/xsx6dU0kwIgdhr8RaHVmxBK
ElOYn3z3wTSh+OTzyJnh81ax71n784Ec2sBWilIIgqVaGbQMpYzmrQDiCZfMApsxqpZHT480ewVZ
o+uimAvNsoK+y+gh9AJDkK/lZj2fPXq7sXPUHFIcLqy2H64RHsmXLU+YBBKLyn8UxDXFVyzLpqeS
rLU/3FJ/RNS8n8qN3MDeagEZJcE1K+22FqmPglMlUksSpNEV6EWxI5/J+po4INFQB5C/iyYZa8n/
t+KiT89QZRl4NJ2GbubmWgad0Ic7H4YY9qMWSO/UPW7CAyJvcbKQ1FlXogRw3ollW/ebKTVWJPSG
20QYcJV5NeyAIbVEN5jzFfPtuIeM2yAojI73qM7LfVYDQ7dduWyOYpt4OlOTxKdK9p2bMdBBLN3o
EKsav2W8Hln7ypznNr0umCE1q4Ok4KG6IyPyDPRxt3dhEdphEDlfiH1z4Oh2zkiAhHX/CGWnmWjs
0SQrtU2X0QmfNfleudjTR5MbFYp4cRExOHrZvPpOuikFJ90ecZSr69e8dqDVH7bFAEwa5SdWgFnK
JPlOOhf4rSC9j7jGF9ZVcXEWEbEadoF1xYTkJqw/ErpPIcvN2BCnk5a4/MCdYTvqru/s5Gx1OYDI
tPPV6gaHI33vHAhODfvgx8VRKC10vGdEnuMljI3XAKUJQBx3Gz7Zg5ojTS8yJvCRZA89xXBRoVaV
kPLaiXLE7Ut8Ypppmzp3SjqNGPDqyn/15stu53gVrGUyxKF43ZPD3A1PxV5j9vdunOxXU72hSpo4
CABv4uYtJhhbthX4AM31evxVELG751CB5xUDZb4l7mSLYboQ0etvY4myGNyEl13BxMUlvtrPioP9
h1Vd4C99PPBos6f7XB1IRZ6vyFPFrUR0c3uNNhwZC6IGHPcWX6diiYu9KIAEO1lIH+P18qRsNgtj
lsBrzg8EXqfhyJF257fAx2jZiW73h3/L2B8GWzMiX2gAkxNEAQ4DrhUaBoSOlbItybXtCwGee5nt
CZuG9YbUQ42vsXgF3s4dEFpkRZ0c9vs6D1jDgeVhzdS3EmTcuLvldp11i1HiymVceVM3EhsL56Jr
DhhEfYe6FtthPo+yUj+kZjAnHGah5S4yGhCXMaTuq9Ia+wQF7W575vDqkppWbJMVATU8xJXhpNHV
lEEHuWKw/fVjb10KnYlcboiEmUhrp0UlX8iMG2mmZRFNPPFPFeqxABxk5hQh354275hwiB559udw
lGGiLcEV0vKnT8pHchoHB6ob3pUGTBLOPzuQkzvQLC1edRfOifQX5mEAaaEuTpRbnDJgpi4BcJYK
GEyCPeKIuuq8lTRYnbx9/zxa1WvsyJNSBRcG6pIUUngSF0A8pmOf3AAdW2BH+BrxkOxcUklRAh2m
neHz6y3Nu5xABqFnShMfWYGmPEVZkPBlYxcW8ZW/zIr2EO41eDFYiQXTIIj9P7gSSXj/P9FFjCcG
hnEoaUTXvn2U7oriAeZYoG3ol2fg4TlcIK2+zkXZir2POKsAP3kurApNii1hpC3uuf59j3ztygmL
7FFqn3kbo7tNAQpjB805WgI8JZyx39l5iicBFiEFtletphR8kIAxkq+VjiM3aK3vf5UVJ/xESe33
4X0Yo6ct4IzwdirLbWjoCnFeAVAvHwzT7vekUUo5uohT4eSa2YoILSO3q3vdJpfXk6nozLjJOdeO
DoWHJ7TzXR0HMN3wIZSz/0ek0/fRQ3mT45ikiG1O1LunIxGW0mAYmE1KpfJirF8jrE7WvZ9azUe2
FeDOeZkMgaGAA3JKW2EUT79esg6rWkNRyHJl0fLhbW9uR8FR4m5XvRAvzbnJX7KvLc9ahKtGROtg
Vt3q7KUOWmZJuP1sOafDLi4V8oGdCtjU1Ujr97uRIbPsZEXIA4ziKXiJ/6ToTETQexhzMNH1Wnp6
uUfDgx2u1O5UGppxMPLPPfioQ9kjO8dlKZ4Cbl5GDo7ALuv6tfzThwhq0qYZUXqa3Cuj9z0EWoCe
pQCWpk8aUtojOmQdqxkMgergGk8W40vRYd5pfN40pSsHvz1beyJOAU/EFMGskHjiCgR+SXWDkTqI
jBF6nlkafUfeClL71MEZZe+BSmoJS/OtmSlrKYycIY5dTp/KngJ/u64lxdY6msGB8Hl0sSwP0Bwq
BNA4fZZoVq2vyDoM8OJHu0lXXlxQKHZ2NvWPEHyvUpqGoksk9wdyNjiSf+hXxk6Y4qaAOuAQMSk2
i+RZg2oignAr7K5w27yoZi/05TWcHpqNuIrOu9J7nyEy4dwnm5mjgy2F5Vrzc7aEES9zh8a9dxBV
Q87zyyQshgoIuGKFuXm4F5JC+q+F+tJhCMzGM/k3a9fH40IlSxWd0IczAbObWKGzaTTk3QNmltA/
EjECAvrZvJnmBdxFphWXjCGXERjS0GMSFLQcnQf09YV70Vw4Z6Emf5BsrSP5G/V8U188ogxBOhLR
gLuRt++MmXDETtCHIhnuAvXWWRjUb3XrQzehAzDSulROPS7PzlE2F/k6iNSsh5P7biJGkL56pVeW
6yVfDzlFf+F4UxNhRuufJ0MwVhBU0eRsCyfcWzdk+oa/DJkd7OVLxmFVxeHxADEz35w25P9ZQ43m
PIm6gI1qt64tMwTCC5m05kyg/oLwnb7TGqma2MHQF+T3rw27WtuTRfszV5Sq7QwOw4KLEBSlnxeI
LumMldpJKTDBVrczeqj2X2VvfPDxe8aS7TUQwoHyi8p8CHLlRahDJD7TzXVq/Gw2TdFtyQC1tK/J
k2HO7XNdc2Kk6pFc5U7KHaipcHMx0HVNGoiT1wIKFv8cK+/Q9gE5oBwzWdptyCs2c+AiGhLM9sQq
aBKnU6WmNdsNHBqJL/kXlq8WGxgAgTIFaYcmozfjOpDFye7KbIsfaEfOPZ/la+B3JL8BhjYav4SO
Hd4LXE3OojbiIMxTzFpEZ/l8JwhDPWNZLbjCAiyq7W5E5v2HSwVu1SQjZU+jWOO/uW4qGxciMabB
f0qTvsrID0l/pJSbr1iJ5dDQzSLc1eZIY3wHPMn8IHtjuphuwRo7NJJdIsQuHoF4LuV76P+quuXr
lqrF+I2vsyqOIdzzI2uK4OTxBxqW2dn09VyT8aAXVrMygfXMmlJ7F55X5koZV7ay8xK8N0az6sm3
MoTeSrxRaPUgdUaevAdahapz/BCAvNyBXUSewsr/FSE+GXSZaQXDINo1aeArLhqfjovxEkLVsCFw
n7MbxRUgzWZJM05rmh3KSTl2iuANmFa1x/WsssW1Mu1ZfECB/Bc5/dJlOpZ3VvpL5QqA5Tek7beg
eDL2aw2c7tl1Q66W+YFrNlRDDK8bDEvO0FQAdH+sgL6j/zfy8P6eeZcp9uzcLOjzn8YbLX8Njt+x
8TxFGG4JEzluI0R2AaxO4SJRttPkVhSLjy/tTTZk/k2BPRgUF0leehGwdoaft2KCnILWfdZVrR6V
4/mt632qsDaPXkBRWuSkFWemF+CbHbnsyL6U3iNxfaW2DcJOdHq9F/9+2G3cNmlcJ5FDYODxVJYf
H8f/EylseU88Vs9Ze/Tq9EjSswixyiNf6mqRW37mwXKuoOlZNmd+MChMBEURB0B+CajQbw085+lC
CRI6n0MbjX/v6CmcSpQbHzR58woxoPl1EtEdOxs54QW/0wXRmoDnb5ZCevG0ACY7mpMGmIH8BMkW
6XtjV2v3Hx18rWqGOb8ub3i8SchLmGjwzerz9vdS+PTWvsl1JUkCG/XWVK06IWXQlzZqWVAKfLJ7
CgNSd/MrYtpn5qQ3j0xB09vwoLGttjMceJiElCdIb5KCPNjDoXp5qzNiu9Pvl8qNjfor7q6u5daD
WOTqFcWR+5cSrFzdjf+N4FBUqwIi/l73wBKLVoziPXsMlRXnsPmp2gADlOxWLCv6Lg3amQGJm0KL
UkAvAq/slld7VtkfDLufNZz1Vk5NGBwcBwQukq3jRaXDs8OPabAHZqk4sBbfEG8LABd5IA3hwb3f
qkyJfb0aVBlNFhBmsO+jEaIi8nmUzpzjB3btQ5fFzqqKJgWIjSqB5jSPSbg54MV8ZtNpKK5OJ3cE
C2qAh1zMzJouKg+03bTUA7l0nOjsKutSLiKz9j5lPAub4RvGBqQNgvILALQRUdMXXD3jidsY2feM
QnGuxWc6FQApGf+Ei724UJDTizfDgGtcQSQuxAcOl42iTsqGxqskNdG6rnniQqWqQiIanpM9L5yX
SXFHCcqHDn8UzI73aEE9UIVYQdFH5SBBsrgL8pdjusaCavUAvimVSz1bi5jepjo9N2ykVyrBKUsn
CvQkJeT9AfRg0UGWGiB+83fBr4dZDF/gKHnaZsWEM9co1rzO1o++dxR0SM1RoXWC1qg2fDREOmbQ
u9w0zmcTMKHfWj5Y6xdgzZ/n6Er+iGZLOjRHpXYz/eD6pyxSmhsp6AxhtlK5fIIswB39OHkIQrVm
JbE/e+VRvXMpSNO7rt08A7lHLeGKEcDXAzr5Sv04udJQjBwE5P+jWAq1hq09HlNYBKKybdS+U7um
jkNau4sxIrFnZ1X/bTQQk2w9jxzjOl0tAbH0jaQQZastZHMFs+C+bd3mU0qhVZEa0omQFTJRFbDZ
/4m1R3fHcsSeFURloQspOjWgOsVDy4g4MiWCK0g7k106NaH0iR1NgWkDMzupHP6I+36HdXqKzmet
8JJWQQE/GX9BUKgzoti1A09llmTHkMyumxQGlf7YFplkDgd3fO9qyMkXOCDuZsd8EEvauz5rFQY5
gBv+Dl+XszMiMrCJ//7iiiJglq6jDsvkG2FQprLujTSeodHd3tq0tvwyEA6T7D2w0C+pXKgqIBUs
MYXststC/t+ZmBiGHrz2ulHOUeKJgE/nRQXp8FbeW+GJh8bZbrSjiZgPGs2Zds5rx7NPotB9yJ+E
YzKM/sJOwfPpU8hCfkUQvfVjktN19NSda2T8toogSCH6waXOz/QxGAKb710A9KlXveQzJ/0xlDlf
LsEy8ZHTaPb3qlY5aJtMB/BLadm5ue1mpm4x2e2J6TE5BZPc4sCnmjB+cfnm8NtKlGZOMS+WNeJ+
FgjgerSo9Gki/CUxHEPaFJ3lXep6pFHmOZlms1VGpRR+thtJia0QZAOkZ2fay746RO8vNbFpFGUC
v8y70tTWSBWWacszIN2dWOBU1hUbnHA4+UFCTpaaKk8BDGfZem0u5aFThagnD9WdqcjxqCAcCSJe
8EmEJcZykCvLjyC6+wNTq9u+npNnDEuUEOXW1SUDFXk93KysqHAW2OJIMNzn8i8l5M7xupzR+HaD
yMz4EsqjAE/DLPbpJeD2yadZY3Z6Nw6ekh9DAY7dqdaohQf6xBxdcovbr1jtN/M/WHNn0iTZ4li3
nZs5B69ZAPSXAX95qzt/wiVDVG908BDIWi1UQggcgT/eyxG+dIxHG3Y4SqgQCItzumTtWulVLADn
5N3aLrBGILdxnXYgYXEpDy8K7DKDhQIGUVpz4m7oL5TZE1FVeo4mTT2hVl59r6YjV1jJ2CEVNqsX
e1K1hOBUm3BFbTY08C/sLz3KC0Wq57vUk8693/hVh93csz3oSlJoDRDokgMQ2VHAI1heeJjpPuia
oAENUIP4pRgvurll0JuM5Gxguv31NdiN4m7/OPGvtAQrF110Usew3Ig7tbMPqSnWaFCOq1V6TZw/
6dxHy4cie3Mwrq+q5Ilb8v/eWwPCPa4ZyEjIVIEunOe/pHxgYRNSr26JF+i9Ew0UpH55L7VWegs1
Ug8rozeXJhSTperPEPPoNOSdVJudN+I+RrzqBFfmaz7hh4gXIVWUXFTDIj3PZMWh6QIBuhK7b1KH
pqiH9tuTlrDJA58yNLB1bP4F4jud3tsySJxJJyQvYBgWvhtfUny1in4OC5/9fHsU75kriHFx8Jdi
omgKqf36vV8Chrotqr/7YTHRyKx73Ub60qFejQB31cnYaA5iS+EkLVkVLFkVDWI9OxWXVN/lTF/M
iYEZs+qKkLfX3UVhwk4E2y3hPDCwc8XWwyUzWhR5JPXCk108UaQEaa6N2rp+O0hVkmp0nXOiBWRc
TIdrv3wzPIkgSnBsjOx+6LXDayImTI8ZWipYitOeyZqXzyAmAAwUYtuv0rO2mojhjUz+vBwjWaQY
oZwUO+AN2r/3ed9Mx3anKNbaG8Fz3PPCUUPKmZSCageBMGKYBDGinFNspPSzLeoMRk5AutoHv9bF
CYy3IbXwcg1as0VFfbNuRMpaprM71gNSwyrwsO8IwnsKRfJ3SGM0fsYH63Ed0CT85obGhP0nF3Ix
jwKRaPiyPOfgpYZ894m1YK1TN9GIInXVyPnq9BtIbo+IfytA70O7pOzOnGao8F5AiRamld275/RL
xNjORXBVJaa308gNTtBQI1/ny4XhPjZ7QHmu/7WNCdnx/C1O1Oalo24omlCVOfynlsvnmvDoa0qJ
in9zMue6lk/qX2ncmIz7TeISU/cbh1HKb95P+3FKgFVPpBwsV/cG+msuTT2d0RHUsYfxx3GBx/3I
DzzzLfKhHdMvG2l6dE15jcBumvJzTT5z1f+/5QkDUDyYS3hUaE4Zi2GAyfml0imITWRfOpv2GSA2
wvWXoiXdBKEcL2w3m5+iorLn9UcPG6wQxQ0Nxsoq4IjzzXBPvQKEbYpfsY4ljq0moniZNqUL/72S
1/yyOhOxoa3WGJD4amNByuvykM3WXXti6KiuhIraDpMo4K0K5KJyQSMdWTfq38vCHphkkbGdeRB5
Pu0+w5tpUFj4wIhJLY3ujpFEgLen/8FqwBghtuEn0Cp/Zt641UY3D5etNA47nq+I2gUtjGpMSo1y
lmE4UxFbm/zuyGF1DiUi5jr/PHit39or5+8aWAlzuUc3ylen+JZqDpERt5YkxFDJre2HuOSMr9E4
qL3C2Xftubx9MJiPTCFdYdMw1/C96JuRuM/ewHaKGV4kTlGmoU2peXlWDGi0wqGBA18Z4nuzotS4
jn+w0RQrBoFBsBke0huocM1b6Qn3pdrdpYY+LsGXEs5wSlmfza5JCcgR+w/k1ngd7CVNz5QLz3LZ
6bg90wghLH/ulIi8gnmApuHmXTtrFI52C+CvGdkGRIUPfS3kOZgn5yD7mdrcnxz63HVTM0QlJgw7
7+RtLUZMoBwrBD8AOgoiMucwQ+J7k8MqSLhyE1M36GDoGObYGzEk1VzkHamDvy9/20hXn5ql8OFo
wY1Zt21p1BnOTOxFXUE6YM3PJVJf3Pz7lHuFo4zeG+pX4rG3eKDd2KhCPAZzRPFe5ycZVYYmrJQh
z47nmnbWfJpliQ9s/OBazWSzLqfzGH//mTdd5KTQNVTCnY++WIn3CjRHdG+aUdUK8XLblBndojxZ
bOmxjVnydkfAaO7DMookx+fnunAJGU6xWaAUwjOIFxxpbG4kLL5IvAIMPSJXiUCZxFu8RixaPt3y
BWJBvjAJflGKxkd7DDruO5+xr//fXBDIcT3LxhA28qdisn7xtL8eg20G/3MSLWq8LBChNFVV9Srp
A8wl6RCSKhe+i35yVa4Ra1dOjhef2uSIVazfHwUAQKWBdf0lTtWDO6rF4tOOzhNhgdqOnmtphflJ
k32CeuDR5abcJ7lu/JNQGjekR/bbuomK/QzDdSsWrIZSr5Nvhrk9645xZQFV29HRYk6acIc1zj7C
byLMvTHYjEy7JN4apviYp8HQy6YGZ7jSRdB+/sCSsL2Cu/XjojFmQQaaEkMayOuoSadMHMQjmEZY
aiWTPDTmq1pHauSxrVM3A1vXDAnTNLpQcL5kKfrMSeM0ZiFJM3hIgP2gDYIZ9UOSIWAQm3SwHiDA
mYcEz09AlNMBZ4TK4H5R9wYQTiGQRQ7btKUw/wUzzwl45CUWc8mwfrmuvPB7ePzVbaeSP8cGsoU5
QIJ82DHQM+qRMYf4k808H8XVY4Ha0eQi+2rxH3dkPEGL/fGlwLrBlV8IArEHqO4RPKPsFaHgxys0
GYYUg3bmfN9Cr05DHIiY7jsL57tzBLS8AgaZXOQJhRSMINdIAOZAM0tYKE2iHAqf5kcy2jk9wTrj
vnutsvUT/g+1ePHspPtp0WwtkiVLiMllGmzcZM8sEtPGXWfTjLkw8MEWxnMOXt5B37chKL51WmY1
PqPMMLUZwG9j9353wc2OdtY9Gtc2lG8yTA/9rIiWIJ2sLS2Jg/iXa661I/o0SJTO+NBikGhceHWI
LBzc3+DOdU3WwJ8AEG0o6QaipEL/zSdvoi1BCriBy+Gx0jGPFquxnIdkhXnxcLzWRAzKofFci7bS
PXp06V6tIvGReuSpYsnldx3BEdoOQ7hz/NeRAF46aEskGAJotSUpdnfvHaRbdju1BGg5b551t0gS
dZG0TEiLhOPFTsZUeaUeZHbzTjfuwSsWR0+cbQnKtFa2pYd/aWA6888vd2c3OGWMn0yG1oautZK9
G2bIC1f08F0mZOBc/PoPdUcI6RClwMqLlNFXScCzANy+OKS0aO8YdRTfOAw2zje/0fyWv4jNolk3
nZeKKj0Mw7BLj74iD+jRkfvf95fUhBfB6TbJStZW3HgN9PH5Sn+x0nYBGkK44HeORYX5+Zj/zu9Y
KPPcUa9kPud64Oy9M5QIltAieTpID6N3KzDsMALUiRivN0wfz4LdunBAR9fs4ABRlER4EySUNp9p
6GB97qGZhuus60hl/+HxIo8jM3Idx2W/obAGuflUi7rETCZT3fpASZsi8UU7zkAuy49uiiGM19JF
Yt/w5d51f/PQMtTCw47xPEZOez1vQ/gD73usdXvgk5PClF8ihFiVT8Pl7dOB/LvZeW3yfdSmmBZL
spms+buT6mUIy+OxWbWOTBTmUovfNAoI9o/Fn/2hJBIoqCCQ9Bwv4q12W8fCV5x8ynT2WX5jVGGB
i+Dhcu3l8e4uo8jrKaGs/iGfS7jSaB0UfhCKw7YUCNKLzh/pmi5aUXX4rJnXUzqCvdLcaHfp7y0J
XqC21CyektuGEstKOIKctH61dSa1Fe0xF8N0Uo18BpnipfDGrm29UGO/+nJm+QYs0j8wUs7spdSR
dpsIuPhNveuhThj+nULc+K8olLlLybKXaG2aUAhuNqI/0GV3KAIfWagCtd6+z2oOB+EGrirViw/G
Pm8hdFVk0F1melh9IX6xjuPQ9FcWCQGsz+fx4C/9OZcyzcEuWT5Du9+NsV3KyGUVfyFhG/Xu5enU
HOQgtwCJXFVQ5BYRBzMAOfAjltzJStcZJjmw/7ylXqnFcFVm/esHT0WVd1r8svV7xEv0pHDoxhOr
VbQyS8fnQdbRthi3yUpMABnJ/rYE5xC1rNkCYWCflconGqMO2JRR9HSOoMACChM+Wow7M8Tced7S
gkDqBdb1kEQWR3krxvkFNbWx7QRGbiKaw/kvb+rF6KeDw3fq7YGztSpycMXpIRu0ENqSB7Lgua2S
cDtuwO/6KyVRb7KwEXZq6me2AG3kL7fX7IoK4KrZpGAI37263pnFBTXuSwAT8l9mbXz7diBUC319
RBIXM0KSkzvmVdvxuSnaxi86XFQGSmGx3ehDpeczihU87+aVX548iVAwFedy/l5P4mcbIyAm4Ezu
HQJ56jTCcM/TpxzfbafjqRNrIVp3+VoEqqe7jPbPhptkKUkGQEuZoBJlQgKkeebirNHLxuxev5oi
+oJJPTiN0pPGxpjqSFBMMYsjn8vbYUBrIcekf4qYtt1zhSxeUhCtBUtS3rTaKnMEv1ALl2PUduqn
HkP92PEQnwk9orAFe71hKEPi/eHxyJTxT+f56zqOIHFXYo538erweY2U9TvFyyMAehsvudibjChW
3eU2ucAsOHUFeYPiWDjra5g2xOZIsQvi1UgeWkIR4WmUocUZRfOZT+8GPA2I1mnDzYmtNAxE+Ufu
sIWWJ92ZYwrjutkHwV7ZKTmt5B9Zs0yBt2sR3aAKW1WH5JPj3HXg5fRZC2xCZjJodBL1R87+lUn4
n1FoLk+BlNcQyTuJGgEfQgx9Td4ezmhM7Hm10YtsJcZkIMmmM0TIHP18JRfSRs5VI4y99BHSnKJu
CHnoJCCJYMwrn3CXRX+AkZslD+L2Bc9GbzUpyNB/rll7WwdW7kIWJ57owq+WTIcgTK3j+DDHMOLK
VbSvMPp+EziJVNt9l6MByZcnrOUJv+FtvEGq2T3QhLgJk1fcCShsyeJZsJ+WUHcPav7jMkLse39F
YgcAP9ieG9FY+CkIjWGmEzwuFkunq1b3Ws+fY6JX8j5rWptZIQhMCA4tPguKDEd2E+cPPka402uE
wEa5tdzBPgb1IWwTYvKdK1a0ba7XBbn6OS5jDjsu6/1FKrZEHprefJTMmJA7Q7fyLXV6r8KU4Siv
IEM9U1SOsuUsqInl27dMAtPOqEWKyK1VoWkgHYvYj3hNKQZ9Cl4sJSvBJdfAsgX7GVc3nEyS8iKI
68xW3pMRuBCSVXSsczHoEpQ2GdcJ8/PC/cf0z9ZpSPL9QBmObBApKvtlnNaiV22AUXDPQ4OJZeRj
eIKFvIAiqcR70HpIWC7oMJiQqE0ZaapIgcCljbs3A2/i8LdlH3S8RKHc338qipw7Bo812Mf34ca3
EehkH2YTBmWqJG/XpCDJFJXLsHO/Udt+VZl2kC/Z0wNHxqVV7ut5+9WLonTpTFP7xNRbdtY5ywuZ
dEID3QhXaLGnl6MOHtNUwHmVmvuep/WAk0Qee9Clo+tdrPdGTNhk3Ry2/4Fb77+XdIYPe0fJJu6k
XQeH9uSif9KTAyV9y4ATuKQQZFxAffYSKagdGQxf/WDXdzkba+sskHl3WQYJqbvtRaTDwBDtoy4D
Bi7RoaCkVFCLIcuAUlxw96DpWwdNEnu/wIEcHDPZhx5q7I+5K72e11++S8sZ/sTooZLIp4e1VAzO
GMQv0Kh1sO+EQBQTp49SVLK95MXT7cjsb+L9DmXHOMVKa8RgWC+0eaWn7ZBxjzxxN/VjPGPtUt1Y
OcAac8uIDiF+1SiQTEt2spTWb1ZKxdECdULjYStZRz7op8uBV1qcbimCnnKOzJJ30cHFUPxR5SpH
fJ4HcHor5lyjBnWpUBJ6L0wfQz9SkAA6nuR74e4pbfKS1OJnfBMT6uF2Fi2M6zypNmYCvbhFlDgm
WJ8vId1D7giK62jaIGnNd3VlTOag2mNn32REb3v+PsDvn2sP5M3G50Td99c2+vd5qjmYosletJHs
izMdt8ifxMaLcJfUGHFyUe46tG1UNZXmRVaL7LE3wzW5kTzuG0W6DEBKYQ0g5CV9jQ+LeFYwvJfl
c4r/VBYMHqJAcN6FjKMldis8C3JJdPVd42T0VFoj2LtoMsgZoZRUPcpCwQXYTMCRPGVG3uqM5z/5
16f1TfRAKJYqQ9d2PG60l4uV6wYJRo35ok6pFjpDzdwuaEV/f+Da9byyA6a8Bj+fvjAA2NQYddC7
KXhoq98h67HXKL2AtwXwEMc4/gVJMD6mAWQXHWT8ceVz8SKnAxiafLhvI9IljZAFHoaNz82eCh7r
2tliCCBBnet2xr0JxxWJksg5wlDe9liI4PhFffpPkTsUqjM4d4qbj8Fr6DlbqYIqMZKKeQdnGxQ3
W9tGoEdrGE3AAwOpRv9UPZzo5DZf+z0+pdX8+IVnkUeaEl7PMLAc+Dao1TTPcbQk5B3wAHtXJoW+
OjCwqLtvJPDrJduAES/HuWryrPSu8ISJYOACo0mLXlM8llry3MD+CKgmuiHejwWN11AH9iyGL+4A
FiJdkmDjCLVkQBTzlGPD04c7FACLYkbrYITLbPijouXzzwJvIB0ioD1x3c8RRAfwH2jBa+lFESIj
onpWYP4jR0bWVgPYm+LSaZ0C9mU22D2FJJkT6k44gCIMZCh1P4ZP8uZuzROuwRF2ggQjuhV7YpYU
jd80/Hzt60XU5pW9ObGqOIsgNI6BlpOb2B/OJQVPthFp0xpUH0D1nQrTEeft7a3Nr5SIrkq0Ce48
we83AzpsWkEEvufLpUMyDkhXk1AufHzAkh43cYFFuiIwk9Pw30KA6WirbXOFdTPcSOdMG9SYvvKc
WgcIH2qRzJyIXo/w9MFLzxY3f+OU5R8tB1EILlKa5LYFhuITS8HE9XAtKiRfr1XX3J7l2h59RrbI
CBw2ISUfp7JibI+VfjWM8nnV3/kGEcSgM9ueewqt5rVdfAEasqcgCY41ssqyl1iLeWd6emL7iBTY
V2fT05luD+qbTBJLvU/dFnluu3Tk8oZn7oTkcmvsUOffPi6mmm+zNN1VOpL6+PipQtgRmC3k2MQS
F9d9aBgf+tTYXeJXIKNYasXeHS2kyBbfVUxiH94ND5Gfq3jtRLFRse0KpTdBDImReIrlz4usliTD
S3dZ9lRk8qBAC9xaY0EsucdnoX6FGnc6oq7Y2OeMXjB8GRGOXLGaQIv8MqJrBFPuTyqYJQD/3/0W
g3ajTQS9NtKxd63NXj8qZnS2xIDJFFpzLYvGuifYMJWhbT8u7xCt9JqSC0v6BDyYz3sNfcZ0aGCD
/RS/QcJA6E9u0wQj+eBQgaKhG4ti8ZrtjvTEcGFsxfv9n+ssirucVxFmlN264qp5ZxVdb3/68Kk4
SzdAE1EoEX3bUPmlv6Lrg2DLy0kEsRWyg4ZYR1KFxOq4wA69ADwtFGFqqYhFzt32IdBujcmsgUp9
roQ2hhtnRXsr5vVnZvLunk2tDEjxLg2ZWFNR+TgSZqo+Vkeg3Ur2etL8pLzaAxhFrL+jKtApUzG0
kclndj9HxK4h5xo20a+y8mSjgPQumdsbq3OrLdZhkC7rWQ4tdNaLiQETWEFSdVgQBXhOUcq9UICZ
xycfyeNbV7qJFwtiqAuThr3QUdjmQk1PeJJnoXB2hqX7rio6PL8MmiaRDN4NRdKOJ6kKeHu4tfy2
xJ2BEu4QfvuWqlgbcojIEf1YdEgUyTT3nDj/fVW4bDiFKCpUC2i/w3D+9I1LEZ/byvIbjkc/aQtA
uDYD+n7d8kYctN4sfjiJk7Evk5IleBq0kda/cGZ6WEqc+pXVECgk7dg54YnsFHVDcA2qojUszOWC
Y/e/sikWt47apl39zS6M58vsAveDUtUVHcZOuzEaYun6ckdBD3snunXBIX7jm9nXoDSpjPHSxcGQ
7P0wWpLkmyADn9NtGS7DUjBul2SHzroRBKGXkrzmLRK7mLqEXXGa2qJS0f+ohSIUUF8bGjJLaaP8
4yqKV5sbSG1UsnOVjINePiHj237+PKjFeaC3+dmE+yAGDssp0GrrXm6FrqWfjKIBculTZ0Y/mcDH
PgXwPHk9JScenL9IZt+VeffyLVkS8e4Xk9VZT2oSNZQlvFelG0V6BWA+GXVNlwUb+82fen5KY9zV
JLJb+S5foBvFKl9DQQJdQi1RCjcS/c9X+fs/dWtHfYb8M4iGO6UO/zoolTybujqFF7Sgo7O781US
EVjPAaGEFJP/YJ87hXbewn7FmB8JvmTCUC60Zmuwhu9PabG7YkNrj/1qkg6FQl0rPw0V2yeIMOQa
iNp1hpYhQGCgjOUGKSJcQ4r0GAdqUrltAGlPn84xz89MbaIyL1pJO9OqyLTFdfR9tOPzI8eRmOQ3
0zaCkwKJEnqugzBcIb8R1KuOqgkJIGR0EOx8hhTr8ZTxXOnzl5FbrWvPi2JPglo7cS0TCB6a2wkr
jg7CbsTAgcAyhLN+9NVIm99d0xLY/4RVn+YBe0Ojnd7JU/Y2TohbVrIGuROk8ES/SXK4tPaoLfhT
usRLTgfpcT0Y4ZaeQ1m2Z9ngF6L4LDqtsmzC/2BosXJq6LowpcgsWPz2VSqBwF3WeQKFJ8SJlBvq
3ryBUejqMKw8L0RCdjT2+SkK6zLjIShHXu1FZifvJHwWscFNIW0hWQTZ00ZMAxleiRxWYunBHh+T
98/qMtI6mPfSJQOLM1grj3mqZibJDz30rJ6yh+2LFHWgmbk+SKW4DtUxduz0t9qRe1MaQXZK5eLS
fKriRoak+OGaq7FMx/5aF3TbzKi8JLrSCwJa6I4Wh7samh1NIkjiUJpvvo0IkNJ35VKUXBMy2n6B
VOHh3gu5zbFuvVKfezKDkpCKT60I6Ur2NBu8ZiD+RwGTulXr0Dxye4pk+TewsosDezNHjaysfjgi
DJwvrHluS150gg3lA/1FbLMZgLLUuBELP5Dv/R7JK3VxUe9QFSRMG4PCYOCjIy/JV8WRapx9x7HH
3NkjR6aZ7tlAkk23thoWbRpGzlQy+Cq4ndg0huAeHCCB7LDEW7k+0m82V2ENs9PFkDt8bqM5CuVK
fprjp5IRvsUPALbYtgVJTuaWb3eZkO8TXQf1dmZfoIA7m6bsEGcT3RwzVVzsO+E88uHENj1NgYIl
uhBx6gmBzpUbh95jaPW5vqMIKShkIetnx0wNjyye9yyk37FLY+7VjqG2cg9lKo2Qy5IXHZcSf92c
Mlockb2tiqje8zll6mTqdnok5H5qybSkPFMDsLGZobukx76yULPhMx/px3q0CPJnggXL0IkeWIgT
rYJdpxcAnAi18xQmzcMCKP8IUwDTCv2fHzN8ZWLnAFleQsQHG+k6dBHwrR4iECyx6+hJBtYuTwcH
4omX8gs2913U8FRKA3alVEqJUPPBB4LujaWqj3WMVGEM2q/iI8QEOOgsd4g0hyPZVl3wMomt3cYx
jxpnayK+XnfDUk1vtBoVlfMt1/3YI3fXEVhMzA2f84jcDman02GWLe2kd03T6b5IjQJhHFMCGakY
CNuq1emcv8pipJjkmf86+DDODp8YGMIEHp1sJsPN60+sOkP37C9EuureJJgvQtCh/IL2Y29gvWQr
nVUd6ZrVKG54pJaGVUfdAZ8SFJBfDmPcZ+oC+d3KM2TY47Sc61Ogc4YqTq7WlnHMiZFck+2E0gSt
2ZSsyGigzA7gaH9bqtCxpRW6CvDIECgi0bo3IWEtA4NvraNpYxAWydL+C39NroihASZngTtR1TrE
bll+4vV0uZu1+5L00R+Wc5GOiqJrnq1qInEwYMZHaGprH6mATYGVOL/8b5i+OyA9k7DALZS8z0ay
7jzgpFLJ0Q/ubKaEpFsmXleZcF7Dpgwlk/oSqOz73QjFZrjNP0KLj0ALmEOwt+agDAFsNXUf5baE
GaCOXhz3I/dvE5bGQ+X3Fexuhpj4ZMc0c1HoIZTysgKxWGfot/Fyt4VRiAq5De2D0nQL1jj11PxF
gUpGVhgqYOt8NTU9YmGd9jzP5AduRFc8YJ01i4M0kkrkwpekUWd1RbBo5/wf/3InLlYO09Dk0ZwX
CQKoo/0I+7FFB8fb1PZAKCgy7n6zck1Sl433yRvPyrFR14gDOvftAq3nCs3zo5SKIFvtAjGcwFnw
fA9rikYY/ScbjcOFg2sOmUPMvjkwEZl3U5QpjzzmvZbhcJigWKzHhSnX6el/p+kvz1TTVl+PVv2h
4aYb3hW/cQc3mQFPUsPajpzgzsHaMipzyYaxJaihEXaesxJxMXjcZx+6eI3adFm23YUnhB5/feP8
zVY14pgk6i7Uewdz9JnczEABqXICJK5WgN1wgJmpk+MlcUpK6EE1Qbh/WV+zYJkznj8hHA0vX/oo
hWvvAA1nXSKe5xXpQpBuy5kyQLjRW8iWfD5FKkXkL8P/Lr+fRySH8TCuWPuZJ645fVAnb/Uk0oKx
CTzhI3pD/CVxuQIhOLl59rPnGv4vhup5U1RgieS/AG8v1n9kJtY/7ybD2smeTlqLnXcPbbxuaYeK
5VDD6AgFJPCj06X9AwCn69I/T1m9rAay9gYhK1MRjZEeHcz8H//aXXB2PJjXPX7AVDiueUSh6dR3
8OagalU0NWDpE1zh758gbhQFORfveVJ24RFXLhPefQwB2PzlfmFHUTvOfFn7BB2MlSvIn+WOrp3O
q6vyv03XurjCduLA/st56oazlpiRILAsWEboUBOXj4KnAr6jhAd1XnFezwnrkrmLDf8fQ/3t42ea
1PZK4B7QJIlCQ2+LE33DiOxw4uRtoTvLyyDz0WJL/wyN2vbVHYAZnKIMpYympI8snvHoxM6O7hym
5bPwLcfwk4WBlSjfZlSOCFsBPOoO4zqnlZKKAsp+83e+LQiTOxiGGHJM5wii8M7TH0rWbiJnSm6C
BGk8FUJcIUtOt7G0ZXO6sFgkS99ui0dbtJpaSDSG7FOToaFrocEG5k2j26ElOY/Oe0MiEqAQ04RH
7alHsgFKzU4fogIxpvVmWog5U3cY7vKTWOQgFZjVA5gp+GLpa74boTLgLy8QxMl9PaNIZgX8Ec4V
EqmOoQ4qeRfkZgVGXo16/Px10cbKva3BcVB/rkC51mK3t0ezFti2IGQ3F+QjdChuZrYmN7kK+3Lz
gqiUl6QDaymMI8JVjVYx8JB351NxXUPDFwee5+DMS1GgzauXABcR8lzwfQx59Q94Pr/sdNwgjlUi
Fs3jlKfnSmeyP6XaGWY5unXnSr6maMoTw47xevB/Rrp6TXN7r/AFpndsjlTO0Em1Y/EK/LY0aHNC
tKAYkiSMAMe8D+Fid/TyZEd36oYRvefME+d+K4Y8A/IJwPclSmGxHNfGjQsOfBzFX4kA/Q7G0aNY
mCNu1jyT8RyhvYNEMWgSdnN5G95sboi82lYsBmbltH6+0o4UW/K08iyYwN2aVBko2pNZiicDi0/g
LjGexH/+vjKFcqW18ozqfpSaFmADERG3qI1Xj7MZbXE4Ncr6kbCzoeJd/eKDjA4fyYjgQwcm8LS5
QIiyfbSWs2EnlQNLfSlmuT+5kzCYILljdwbPDDH+oncvO4jvU9BOdSOMeN2+fPk6r+lsMcOkPzYL
TUTAKq/bVZMGnxQtIecdYe45rpUCNrMJVOGdVxg7rbFFhSrgAGmTgFg5pwgPLPLHWV6LdP0hFcFK
mVKXNl+FLjXUjWYsdTY9O1P8z8ZKrrc1XfuYD2cEVYT97afM342TC3CAAc5jSlWrQaiuL1I8P1R6
+wzhOw9ajBYEjbfTuiyDy2gjISxv7K2UbqIt0t5+HimbeqOuT8YhSXFL409F7u1flGj3R/Gjieqc
a+69VikfCW/mrVwVbej4OZPTUfstuefAHtyLZ1J/mal6UTIBM4pEVoDna58pU5uY8pyGEMbFlmQ+
KLw0S2Bqw5Nb3YbS7BF7dzx9XihpQHsdYjR7IWUx7sK8xI6S11IzGvD3ea1vBSfQeiMwx9we/a7K
P8u8c7tiH1cllOTKv7bQW5IjDbSrza/cDEFEBOuZx26nNxMMuK0JEi8a4KRlzcdYCwmSZDttSiXx
w5Oct29b6Nu442xwpIZrNc0EzBFjyGYbaJuDdGBBEkG9oAhgGFWioYI8sLV8S1jtcZwZ3oKlbXfc
X1AqH6CgmsEkobn0A769ZooT7Q2f5wNksUjjClo7+DkzM5LqJGNVqYleS0G4LJ6bwUWCrKTYTEvR
ou8XVFBAl5o7rDJXrmrzYg0/+Ba+3UV6Qt1nAc6jUugbfkNYFyoey7BgTjqdL7/iTn+3M/xIYd+W
12VLe6fd5QgzsbqOSGp4WJ6zP0H9QscePdDIZuI4Qt5RaaUgZu5VvAPmtjmDD02GRwq1dDxGp8wd
ZUS9rBTjeGxRSgOQUYplzi/R5N+FBoPOlVgOKt/vw7PE/yzIqgA/WvxMO3LpShBOdnG3pNjBt91O
cbKPczkQcr5IzGE9Mrj6YLu7qwPo2crZzvnlljCr9z7B2+V1vZLnNPTIysCcrmLP/Q6XV8gtS7ZR
scgAe3dTyHRDS14OUOTHDvGQrRgZXzt/EPMDBbRHMwGuI4HdARvYf6/orQP+dimgGk2HY81uSt91
NRLoUAEc5cAKNiXQSncE/ig9mL/3+QOtqsHlWtFWgYxLH4S1guZcbvq7MW+JLvK2HSmd4JbHk7jy
ha1eW7V7OsbCkKBixJrhiRpvIDByKyLsOCHDRIYDUCxpZlyXV+I83f4yJYGO69E5ZugmGuwzmmWF
nZbBmNngbvsxaCuYTY8WY5GGAuQ+VO5V2cPv5sGdJ3WBxXD16eUHFWdIhS5qCVWXSPWNxh4prz9d
itGz2VA19Gm1CGaIrssNRBvZBY9FT8uN7q9FKxvzeYXN9N1eTKgKqRlq6nwdatxJTBcUuvJcbxuV
UVrEISroO+nKFSF6jcn+nVRoxl0XHeQPW/WZvFNOsHSV2Y5wa9VhbeU17DVI27XEybNvj+KQrePA
TcuMNkMAqY9sfsP7j1W9yXhbtPEu1HOb9D/BDOH3YpAQK2omusS/CsnIM0tsFLdW1TY2H5mFeohk
CpLmJRDLAgX+OKpvp8Mpa2HdEfq0rFN1WUrw8gbEBQ/Z6xnoU5WbgkrOpiYviSveOIUXarL3bJRp
kSS06KvLQVP6ZhFk04f6nhxdhDs+4k7zE1JawwOMDlKmljoJOt7CgcIlndIynxcKWYovevqdRj48
k70bhIK1w2he2AvtWHyVyRIVjM9oW4dHhrpW0g0AR8f4nVdgqj8ENtZ0BWr+k1OpG6vfzHC6aMKr
EDfaaeMYRJk4ppqSTUY3QcofVo2AuR1GOraCvogErD5wx7NBSBW/euBzx1QjGagOXo9CweFWI6Wy
7ytmVYy7XOygDPc1hPduoiHWDjlnXPF0FKI4DIr7Jl1uzU41rci9GsJQWFpi5GFVzZBt+xbUtsKV
CTEdltcMsdbLlJUDxNVUyQMeYcJ9Z40HvKRgzkvk56nezB+EdkdEtu3nqvqfMMPDvBxnS1WxkaZv
g5+0i1psUzgxlHDTyqcURwuLDkyg3SBNvt1EcWqN6y2++ZOWv/LZy3o2pMcs1a7twaslW7S4YqL2
Z2Is6SaS80eU6+yZuHi7fMex58xFFTSamcrBikXdfQCkoFjXJSVwHEea01PNFnLEpaig6RKA8o9m
StiKRwTHC7goXp6wM5cC8G2Mn1zpCazJiqdX3ChiuUVIm0/AeYMD4WgzwMIG/w7tRjnH6bV/oAjn
8AV0CRE6V3a39yDTMPPLgM34qO/PD72a8yc9J7Fs5MMRypfaS5C50Nqgty6pPptN7DOT0Om4T0CL
xExr0nuHOrIbieFLTBSG6OM/4bff9v60YWzj3QE8GFMeyRM8WQ1rnvcoRC/DtF2qadN7uZlh/iWn
BEdAV2maJ9Qj/X4CcqdOGsMQeGWaXku0mnZCbjR3jF36EuyerPMuM9wbiiZyGBepoquNF8EX3jX+
E/PkPkRSWqiwrFFmfM+5L3SZ6uTCQrc7Opd31xBf9xV+pezBIQldm7fXNiqe/X6CjBgnp9vXECUW
ICLR1o80Vu+H3sQpJ9u8Fu+VlfH33pl2NVHWQ+c7EzfPrzvofzWLawiatfmOsuTYrPJ6pTlpwEKE
drDtTDeLsx7NLjhPim6+Y6Lc5EmRO4YdtsK7K/EQQ/OGVPPKH+E/OW7Xu1drddYFLgw7pQBGKvJz
FYd1HIVVU40/PAA4GS8Mw2/aYR/1kN9vcAoUEMu3S5RVqiITeVhR/mquhUG5oUHmoRvxyrny/lAg
xM7qleABY1vEZsrzAIUqLF8yyBfQMEl5CRaZ5Q74Wl1Wf7SNvFtH1AK1tsvLoP8pbYDIOeg/xeKK
80YpzJQTCUnTYsj0b/zE5lLLw3OAhajsD07S/AgWLLPsSZl7o6cpUCFSJQkBQIUizcwonUlGIavP
WmL0kR/Y5J7ZFLoMBh1FQ9k3dt5krkEQKRqS/E8ZbTGe/hv9pgzEqQ9ti5po6+EzIHG/BXLC1Hms
Crpn5DsoRsPVKl0R915P1vXAbF+xqBp8B8iHnTgtk5yQhBN8cAsZXA+B+aAkEeu27JoWPKufx433
rFdBPzYaeK+kscAjjZkgFZPDqaotQ8N7w5F9EPRIey86qDRkX+tkjl2KGQVLFcBCuGq4/L3gDovA
jWOpAOhP0CDAHmwHeEF8CDwvWPXULh15YcLedvrzdXDJTs8dFTb3DYGkKmO57PW75d/z/+K3lY2O
Vbpu58wQhncK7R5+IIlcVsWbTaMjiZ6/F4qIxR8LTEyxLoAfB9VeN/b+FQr3D0sxxSxG030g3JEv
AZs3rklq+So1nJhs88Ap0LBIHzqwPwVQrDzu5HDO+XgsUGXcqZ9/ckcAiChpKMCrtCn46c7ibH+e
CA2a3VrjrGzTjmIjooC/buf6rMxYmzHj6Y/DFscxwaYVoeVe6PnO+NznhaDw+o+rXt9jsXmJQ0LF
1DhWHMFhwc/BZgihwJTbNnL8/CAqGWe95LORHvX1e9xmNYpPJtCQwd3qP8mMrwYSSlDUFAVrKwpG
XLjWlo6u0SkZCOCv+hf3LQ16zWqqHC3/tTxeE3DTMqzyMttjJU90Hz+mPin73khs5Dp8seKo/vpt
JN7S5O+P7gVY4ZRg8mo9TC2GTqaAZLO+sTW9+2e5FLM0m69/B9dyKOgBmxezZhra7Eq0KNzCTenl
V0CcwmMlKgh+es+e0oFu+pT09M1iw2yhMeyP98igDGfRkRo/5Ae/a8EEX0u+coKFTr/xnsk5pfRx
zH0O9izZWx3th+rV2OXbOXQdwbPS//D3ZeoFEmCT2MLrUQ7R2vQxNHeM07Bpy5VJkzraY7396JCn
ZQCopkdSifLbWIBK4swozdogDb8CZFjVLKAUMju9qZSdVQmwkP9wtDW/vbLF51oPKj07FwwsflfE
Qm15UL8qR2R+ow6ety2enEWm72L+QzVB3Qd7/06qsRe5ERBt/SQ4h+OuZNnd9OdpML6qQgZ9wWKH
mHItMlIpJetcMkQdp+Pn0nDW4fiQ9t+ysYNybL4F5myhJyoE9dTZ+PYtAWgviEcDA7lE2aRyMMby
bnxyFFqDyvQQ90YgODBGPZlTq6jZ+3Ft/syhs7I0Ht2iVNTJqEJ0xSLFya/5Y+Mr2k3PusTlBe9I
//h+oMpxIFq/2edcphzeg8+0UDZX1usbuVJR7IPyuh5qOFz/NRW8FNbKK2sCTV35e9rsL02Gi4gP
N4f/OEC3+YVs1hSBpnncGsoS3koTblOiL3UN2qvBPo9DPVp/yKXOVX+SLbL8Ze2DfiE2ik2NrEH1
g/Glk4HB3zTiky3/780OxVFP0q4Bw5HVp3K0vKaT+tw68QxQrIwQaHfnuo6TRAObAbTD7rKPIoUa
hqL3jIe1NHxR0PLj4VOtJqyQgs62NYlODK9MPoGrBmXfGjYdDFat5gbNh9U/yRZpeUuNOn1SHRoO
N5cZ7TpLp5cnD1I5o2IS9vY6gDuGNN1SkMzfvBohDsTsUrH/aJujXW42z+1blP4dImgno+72SzJR
gYkf3xsM8jz/fcf1hVWvDqXCMAIVMwFqTRUVljQLsIJU5+cj88kikbdgV9oiDThBoA29gLfP6TxG
u/yJ9poKw+ETf3oDHaVHn6woB4ajmFXC9PwxwQX56SsZUQM55cTl+j+3B8f2KjpIe9EYerFGaqV0
p7BlOpBRPHV+Ucz+NdQsP3ZriEYgqexR3NcYz8X0yrfD/ggAp560ruM1pW34kxQkUDaTjMvqM0Nl
7wl8iJPwfVAMsJcKmLOroRXSzH5hdfRxemg2/oyJKgj8J4ntj0wO30yyiTpymmWPLSpcXxVJQWL4
s4Ownf06W/uFLDhwYE64ZxzynrNgSMhm+0uUspWLUdrxXiUqM1bulWsyOQoq038TDk1SzGZslX1C
HzLJmoP8Krj3Occ8Ns4DewCwfVgpOLcu41eTQLJb7Lu3nyTzHnNWStPIG9vtc+umJf6hbsEbY7ab
OTej4rJ9ZPY72XWs1B/Wpwa3PKwYAlSWRncHOYiHb+jgynYJsp/DUJTuFhxHNYeowTOBjymFV6As
k3DNoF/CY8BaEMqWU4XkGOUmnuNox8dxo7zvhQc8cPrVzhagav6UkzWzT1Wsk3yUWRBfP9A8Vw09
CsQlX9sGfQLuVyRzMOf2yb/46sU1rA481CbWoHdxFKUmv6qR15PPx9hUPRKphIysU6VkPK4f35mo
Mf9FHyrgGkF7mK1G8DExhdLGog7/fm7e282mROquFI2z2c3ve2Pf9fwtf9UUmR4Mc3JCBfacq1M3
6UDmfvf7f2KAT83fXEvNRlwWIi0GmJi6FaALP+Kk5h0b+iuDek52MUZKNS8osItapbk7wz/NE4vr
jNhUVpOQh+4/lVSSkIbkum9/xpGjGKRh6EU7QKzyaYpjI/dd5rH8EyWNzVQrvUauik8XdcjPJsjS
YPzPpnsuy3pllEp/90WfHWpXBVsbCuCrDXZU0ZPBotcYAT7q5qIZsP1dTRYWb+nix4h4KEL9r9Eo
kdIdt7owVgLTG+nm0AfZkx/aVEkd+nBUxVBq4aUOEcc7rfajehqy5JSOtOLvpBAPQoxv/rbVk6iy
gnR03739BPQ7BWZilfjDooohdsGs+HUL9frJSCXMLABjCz06qOE+V7EYQr9O6g6B9dKAQ4N/MizG
S+qf4SUL/3jQSG4JFyHDShfC6QZ18sLjhcs06yZNLLkVKEwzPUJps7CkFVeE6StpKtK/Y0WEIpTU
P+CbaUGYH7nLoWItC0SwSnWKvphQmjnH6AOqSMhVTsOPAxIiI5Q4LdzVmg46D0t7AQilDtv6IScW
09F2u2gbO7aP59AMwipfpOnn1mpr33aTASHbzbGqI1Pp9K0m73Hx8hOQfkDigHU23nSSPN44FLS0
JNlRj0fcZUj+wlM1fnZ0ceomhcBLLu2vrrfn37SttNLI/8h4dvd+VHs6F2EtHIzb2OaE2gQqKKhr
ykfr3GSpxozHVBYPGNMOdpxRmXhlPgvUtreANLq95x2+9b9JsxRrX4Ox4bpsIOuqUnQPiE+b/HtA
2PVbkx9k7mmlZo4ck0c+Zd7MBDsu1DHMqcqJNhMfeyZ8sed2IsCuw8/q9k4+OS8ZX8VjwmZ6INHh
m6IRyntyhLkbnORw4wUpydOXmlpquf+vpG3DPIsta/wYsJcXbovVXPGQLGcUUs+13TcZEsjku+kA
rcoJ+b0FGcuYfdhUHNJmUkL/y3FNAnBS3KCx2pCTAJwHI/KOZNqIQVJLK0d81JM4h4YuSoY2xNwo
SmlzhRSpdGhdsyGxGp8TIsS4oJA1nflh/pO+xdFMk7kvMSRsz43fs2BHhveyWdrSspCVmLgH2B2Q
PTiSQYaQ8+XoYZiPN2/lr1VWswv311YRvCIKIpINYfxTUMJ0wkCsTIYR9fK1WxguXQE9iyc/h14D
64Ti6Jv9rZ17/o4WTh45KM4HF1AASoXKqd8RjtLELjd20KbmLavJqeepKNFCzr/NqcOn/sl4y9cW
zc17DLW8XzokJxaBGzVwe9qImnyzp18VtBkE7WhufQkH7H9MKbe3zgq69Dhppw2SvGsMobTM3ws+
F2l6NY+cdXz1nLownHO7BzFs+/WjPxUWVXtX14coZog9P6Y2WhiG5/A4uSDGjAQS7ePNNXCAM2ri
CXRtyVtcGx+uXRGJETuW5R9Pzx8hQyfdOmv5ppHf7LRAys+Q+IvBj6uuYcmEKDW5HRQk08BMK/KF
9C1b52Fb4r9PUSrImd6acLzW0A/8LCCi4gjuNkzxYj5otvyETN2DOddx7Zts/qqYXWH1qxAFxAAj
Tz3KZdt7qp/F5D5YSSWKnxCnePl9/uFUlHpK4yZz6IHhjLeaOiMwJgqqQpdF8OaKOgxEEb84RlOD
LFAFC51DfS043fM0Ff+ScVnafbVOIAXjhqBL39apLi42tJzX9H0HxmigaNrSMR5zFgVlVCThJROg
vzRrJpWQAOzCTYYyq9dhg3bh2DB3zGBGNTIDW7yw6kWoB2RT+8shSmvJTp9Zhb5Pre8VcGvJgSPQ
nnkaHHjM64QyUl+8cL0t4jf/FiNyKTA49+CmMY9RpBk6RZAxLexj16A7ExlqZ9C+M1VYwLzk8ZF8
s2c0tJpQ53ZiugIfvhukbxLqklsoYI32x4wOXYbMOcDc/DhfEauz6jdguhgSJxdB2m3qikpn2Slr
38PR0uuNY+cAJLw9cAXGvdnfQJXA85/J82u4uwG7QH9h5aEggl401H3HltzIBMOTy3741mSEaX19
CAX8fRtucbxASjlKluR8whTBWqRLqYx607BIrXxWG+7kf+q6kwHk6fbSFJCns6uc0P68ICk07pbW
tLvLGli2SvfARSvBK+7FIwglonNCGKdNl0seQMziAI8gfn0iquVFaAhjV0jdfUIIBwlDaLiivJaC
3F2JxeGGfN4AHL3QW6O8dX7q+IchTsQ8txHghbQpW6NEHiKg4GSGT+009ZhP/3Cl+5HaSQ1LejUT
7msz6KhmXeE2h0rvH6hu38EfGAa2MfomKWS4eky1g4ifCxd/HciOwwT9dWkx2zd408iTW72/K6Dd
qZMPYM8qiMu1iJ+mWc1DAb82Z73BvHloSWZ1uAif3+3hzcLIm9YbL8bEyKTubADb0yoYwchdOeSy
rgbnQscVi4rUlqRWCCvEJXMUbU2eT+KaG0VqyKu8rPXfKQQgFLIgJnMUT0wCZ9kdDsTulHRHqPwe
/3hkG6z9uarS5ZHdde2wsiu3yovQI+f1QXICdhG4AKZ7aM63QMQr0ViFP5j1FvYZcTKxCgU4Hm17
KfAvYx2u9zkrqZT0X+nBNdOhuZnPi+rzRtRbGT+drx8cSIaU1g97II0NWasG5+V7lsNdGKi0YHpK
1MhAD0UmVuCwZAYoq38lwV+SjVz00AyB4N/52I8y9+2EEEKpnoXRJDc7q3V1dMiXi35+PGrwBVqN
DVHjk6xILNsWi4uuY3SkAWIFIrDTTwec2csFDuf9xdx5ti5KQzfje8fOH2Wx7vo8WqeqGKJxX5pk
nGORX29eSJBaS9bz5LiQ59iWIC7YdHfLR5K5i1KxEHXgyPYFbbx24Ppo+j/tMRVwU+cuWCejS8+x
vLXPIMSyKX4ZiB66zrqH9QMwBrJiraalGnzsUHKp0A+scaqpwCWvFQiHCm7XPm5OGrC/DnVk6LMZ
4lrvoXlJQze+iuJCLMdG9L1BegJsvL0XFox/KnwjS6Sb1wPEaj1s+A6/kfnqSZhn9g4AVYLVZUZY
mjRH6wmiXYTWeZ+Fk4R/CrCOcQw5V7jxMMnW4eXw2h75SSaENJXh2YcBdai5epZRAZnbtXhKVzIi
RgybB07Rqdf+HXEDn1J7lcladmFil1kaPiVIRB7H337+ugEoREN9nrIj7lv0ik0lLerSrtK2/NE7
QGmITYonLHc2S2RcXMYmX4W2fCRH33yg/M0IcU87eZtksdarATtvsqJ5smpVQXJJIleP09VmUWA/
BuM2VdltyPL0JNHfGVFCJIJXCP16G3lkeW/qeOcg3B+6vn+7UQK2aAaRbEsWzQ4F7Ewa0FIQE1HQ
97u2DkqqjLrcMTJEZHEwggV4JuUElL3hR+7ymtUFACFaw2kh4ztIWW4FpwhQ0Y/agB6WuUgCco2o
SzKjYMkzToyJzYRMC91xZaepaeHp/UttsYtgSPc/NzWGMDdv2WWv62opsvnv74nxw5N93cddc1Bt
6woiaxaSBX8HOh1/JTrWtk+L7YaZfhpcjKKggz3LqHAyIM3+XQyhMiMn0Y9mtfxA0GC8GDdzH+B+
rktuLtGq4eNzdpcmWHWhBosfqFb7V9DEtYWYxMusfcwUHh3anyW5afwQC0QuMLUC9h8oQLiNNt5E
W0lB5gB8KLS9ct8VcxAOQWtfdwwHeoMOuEzqGLMT2Jm5yreZ0mew2LVp1urUuRSDxPAXrP8Iog7p
gm9vTHKcxmpFPsxcLQel/G0cG98loxBYiWeu4IgLuyPDJn+wUV/ijbiCa8nG8uOz9u8sYAwnZKN2
0n/zLqyfiB0e8uyOysiyh1YLVQ2wY8/fWVsjmNFCe4p4BndsjcBsBwWDZ3O2CJPT5ZUTLZuZllQG
XZL5Y2Y62CWnZQiS7jSrujlah87Y19Zrdy59ioeX0LlAWP3YQs+J1xyTuASXvrIAuNR3RSyQX3Zb
/vm8YhaOEDP5GmSZVyVbZmye2CsHTJpHDeYDVVMpjSei3bK/K6yUPTtvnpxYPEQc4E4WUwr81vTt
jByJgVg5fWtSEzJyG5pAu1ZZMRyBmqaX8AYVOGPtjCO+l/gxvt+gQhuAILCfYvcQ1LpJ6d7RCtzL
865nOinX8umeT2X7wcHhrLosNUupf443EfK43webJLf2gMy81Jkchiu8idtyL7prHjV3HbUUBVsx
W4okvmfDe6lvNSZ3VXP9y62hbIULqyRAkofY34bB2hhhHBNUDoXrHc+aqFwCn9i5J6R3ZxC1FpZS
8HCTZhh1rymObCOLgG9R/qGKfdiw9PlhbPpKCQgWECYXye5DDSHQ2hZPRPGx2aaiK+bzHHeXvwHX
7bks0J4Ys4F77b8Uc0PMXIcsYE4vbWKdH4Kg4h/6sahikh12jM7YJ6twRvjAc3OHEL4s6MnjplOK
708gGEX2BmIKtnin23YcPxVIj7uQRhskm8XREBoVyh1YA+qJ9d8ifuFxBxzkMBiaY0Hyt2uxToYB
rrl686h5r8/o6PjtJZPdjQ5/2W9f0Vlhn1O36gAJN1pnpYRZ060q2vRMFkH9pNxRdAD7kGUnvTVv
T1b5kiBgHzqpwLoWkLhx0L1Ukq1TyvJI4RyEAqw88vmgMfJygy8WZYA0bijWCBv9O12dlf4tPsgh
w70Np/kgApZfkR+DOxnN+88afFPhjl56O3CNwMl7hOn09amD+kmJW75Avf7zZ+Gn2aqmrLFPwAb7
K9h/IzPfGHV6LEjYIG4+YxhwSAv9ozbrQPlrL4y8TKw8q4PP8qZAAUWtIOjA6KuoAVBkN9GFAJSJ
Ot/25Cj4mlXVKJuUzNG/7l8KViJwEO552HuPHeHxqiYg2b81akqkBPFcgRWqVjBMfBv1OrpHHSMW
4xfiLaPXPuQnUaP38hE0e9SA9Q2yYV1EvoPy+bDBKQtFL4D3fgCPvSQaPGg/ZLFQY7ATVtHrrJ/U
UVxJ5IKGMeO5mxtoKGqkKumCL9GrxJL35rQtl3JEd8GIzjZYLYmC76Eb4aZ+RjDhlDzu+c5/DJka
nKkpHYxM1uZ0uI368UIHuECiNWRSp1gKXaCI7ol2rngFrMV8f6opboGVMTCDsTyfH1ut42oqqrn2
GztT69oslymGp7Afl0ZSYxRS7/jnRYTLaExcXX1cfygCKu2t5OcwL1DYzvUcdwsqBk9ru9ixOSl6
xf41UonZNDAnwx1bX41aSK+8L1C/3M0vxktAfFbd9NxGCgz663ulXeQgePWNOHdNJ1f0bADrQPVE
8VPXlDPfhqGxaZw8pIiJPlH/S1SPbjIezjoGsVFs6xQHqGbFaYDIK4++k7FJCaSSp8DPrp1rTRwR
sV3/y1cQQBnGWdNWiKParDnUfd198TGi5zs1ZqY5ofsiTHJjsa1DlWR6tQDU/rb7+cYP2Iiltteh
d+YrywIKyIjO+2XtnIQgUPfhh6aX9offQq86M2NYtQp5nSTNOmi3WPVCJIUexky+pjlXg5FoPFGm
Ccvm/shiUzx9BScWfP3Me98DJrbXiQJc7Jppi98PSq9XGNvJJ8rDwjBOejFSwps7Z68E7y/YHRDp
Wv44mNj8a6uWuYdGHZrFG3ZTI2XI8tDbLTZHfzpmkBtEktZ5Ns3wlCtdLYM9tNElZRMu00JO99iE
T2H+NxN4eeLzKVnVwN3N8kYWAOobfC4aT0NBLCtstELBhQZ7AYa6A/gKC45uPl9p3jZ426NJAfP3
rUlWfov1pnezkT/koyR6J9PdgIm2tKLb4yw/uHCKPebN0zxx/glJBYnsZ0eJv8XGLOEhsWj8iM0+
RWOQFGveCtniCmqJLTOMpvHQUDPgCQRw1lJSV6PPivvDuvexwOE/tP9ceRnOAY/Tyc/q2PnrBNZv
Oq3+87p+Zyuns0D0aGEPXPXS483B1wRauohy8l8J0RyB/UPt6rVPCCiRAfWzofEFfxEy+ZcuquJB
ylBPAJR4aLenFaVctDzTanSD6m+r2LM4qqmuosHofkuL6B/DZ4U97LbvAK0szlCA6sGbpyVnpk0E
36n5jEDouX9AyBQ3Qh39ESM60U2HGg0mi8cVQVXBJEeyJB+9NX/Mu4H4OPceZIuQJJ5MzV6g2kn/
b4F3byTebirToiGoE6acRVSWbYgYE+cvpRAbhA5D208f16OZWxcVdWKU29bTSyzhkYWw7doHwC1V
ugM+GphyVUSA1u8QWXvxVp+3O6fzOGrpwikIS5YeuaMDc7xoIxemQNMaNuzzeqAlZX9hAc41OMfQ
062w67uea3b3A8DmQunlZeDFBXDjEQL86QSRyci7YAW9WGbVLEf9W5KQP4cuPX2Lsy9IZZXxNFUi
6bsC3kIF0HGAGygkyA7oslofa9MskTWbTTXjsxDZqXAnPno5lVu6O4bblWwHmOVpvQUFxHAT11IE
Sa4LTrXKq+5//BQEIcTbJehTtdUD+I4YDpi74UHVM5hS1EyEGEt7Dmj6TdRsoJwt1xY0iKmVRIOj
sa9/pYcHlkj2YkCMkH3dLKKUu8M5jGwiW2IagW2Ghu9cFssyE/yO+g4jbcfxzKEiQ+HQXQH+W5HU
MoaoVwg9AK2AntIuwfB0vP+oyBdUGTInZmWJNaofThZ83+IAR5KWsG8228gYmXt6d5QqWSBZAIZf
MYpXZRMG0k2DgEC7LfecXDPEp5MrxLMpu0Fcb0naH9oI8YjEOPq2Yjiq+BQwdzQ+I1PA6UwA72aV
3Xras4Xq3A6tKlfHCWpEx8B+HPX7+tQw61Hjmpm18MNidjSfstY2lRPEiEcxTy7O9ceSvlll5Ykm
XYkdAqx5jthFoSk5Ihpk1tD7sS8yPR1AGj6k8IwsUZxZdt1MP54zePMN8M2Ri4e/chgHjhLNFFTN
1lvg4qvG+iDOJk8z8WfvboQaQKe3DQdZZLq9si1L5whqF9pC4GHp2d+EYV80Vn3uCwltnJFYOy82
XZDyP95PTsYXR07zhL5gv0Wz6/e6jgiMawPPlFY1m5Hn0gzV7+7BjKpm1xdjBWnPWjiCBsa6Xbaf
mo9vqToogSVvb1M4torPKuxYiVcJj4GSwWJzCvEnka/vUJ6LwGJTGRAS7h0KgMXut8sHXMvyRLSQ
2G8xApaAOrM+0Li2C6Sepg6r1RaNbZfSH1SBudbc/nY76q2n5rbEwKtENHQWh+JYAFJZ3xZhemt9
geLeeoigf1FSdjfcNsj9rKIZpDohe2pWqRBY/2in91Kepd8vNq+29++W+FwP+OwhHPib5DSQSb35
MPS5kxs5V5pW9pIrQKj1YO4lhLbn2M3pJW5UrE2wlVhtE//6B0QO+MTVQz/KG8KXAl59qZnGaLpA
Gfd0JNydrUMtbMyM/vmFTv2gMUSf5m0ScVD4k4zngDB/x5ib/k4H9H8UjSUrj9vT5bmj5WQ+37Tc
uyT4lfiDj2OZotLH9T1Plo8MAUHt/X17B1cggqeaF3Pjpx8/LJr55M+5Ij1/sB+JpZvx5Xl91Qqa
2FNqlFvywYA6hkUKODWqGyZZ/c3mQsBBU/r1RomEy/cJEMZL6hXAtqr67ll4i5sPBFDOmXw1m8qp
2BhssJ/JkhucD2qNDO0FJWjeWW3LXZqNuYv4mHs452ls0qinJllXsuK0h9UbeN79x7F4xOR7Cxiw
S5z7wrurSaSB8gOmlolFhpvYQ2iXUudG/ALKraCJqb6YOsIcd4dCboYzz1KhBTqr3vdw56zS5zdr
hRfPslgLDVGoBgbg/MZbWfvew/JMlwRZrzZhfu2yEnN6j1tsxwa4O2z3xHewgMePVsEKOjF7w6ZL
hKtV8rSMfem5/i5NHyCJCzYxap9sfENsfjRFHYNyTrIeolFG9ofl1nrETZ3VMh3v8SkWNTcQUppb
SVASMX0mUO12AmrvRbAC2B91abJ6MzRkM3CDDt5/0dHKCBDOmYQBB5KEOy3NXc/9AGgc5S/KezV4
arbhh+trSiGsf8ZoF7Tt/3//U2eCGWo9o60IoELt+Hv/lG65XQYuvOR4M0siBFD8m5D1xRETLYor
sGT0H+1CA8HfMTchmRj4s2Kny83DhW71WBLg8KWvpb9kT8afnr+5UQnd7AuZNDSWLrqgBvKAB+00
0DT2MN16XZOWJuVM55sqU/8XLT7tj4Ni7O7X3U9RwN5nUS9zs2Kj0NPesjPo+9BRgZeyERp0Nr3S
rmNeSIACsg/UtZbF2XXISht0oVKm5NUQEJAIjkUzKvcnkhHYwg0PhFYCXtSrgD7wgBRXr3MTcJ+Y
eKzi7ZZ3VfzsnfoGAWJUZaq7/fmT37BdcT9bUBH5r9wt5xdga6AAN7I56HiHKT4I2WI18/Fd3kRe
Duy7VHNGKEdX6SE595eRyRiBLJkv6uPPPsuAfyZblsONne10qbhXTjsQ3xsBTLcTHo7Gf7BOSXFX
CsWDhPsCzJTgMMkaKd6jYhU0eJ1tpEBi/niavVjWce7oPXfco8moktgZwKIUxBiV+EdKUZwAZbUS
LpUtAAuiSuBwpo5dnUaoqOMVPLWOa24O1owSI3xc1tx/82yNROoKNIb29VsJOYiWVtqioUp/HvtW
+TSe8kV0KOCjTJk8nztViacc+YAktEQMaumCt9AygaTf8cFL78twyiVGEq9y4BMdIamUSNKSnUOg
VjLUcz+hsVoaNELDL1VHAI1EFMKl8IvNvdj29uZPGJouP7crgL7FYXVIagLp7ZKxp789elkW84QE
sEZLI6RD91M0jU5ingvOg8sCV5vt1TG2aSl762IfQVprz7FcVdYppflEd/Db3kItTvXjeVsTnopP
+7xzIo5Vz6+/S3X01AU1wry8HRgPORO4AsTgCCPeWy90J/AORRQn8V6yddfOSN1AfFBAaBR1WlcU
fmNhJBSpmyQjW2INl7hxOTqMU7lc8q5WNQzME77LlvqJdQ87yzjOlTn9WqBcc7/cnmiHlaO9gCbH
RzUx8vsLZPI6IBjAaz24TZB57CQjeyZHRathGF3miMq+y+LC5oaD2UKb6eOWUnNyhCIApkvNLd11
NiIR111mqgpeieJo2wmZRYtlDxuBatWUA040Ya7i9XLnvHt2gkLUWbDzNOc6sQsOgKvruZYnKXck
YiCVyYHAN71NyOVg7IJZoy+vUn1P5sEZ1pK7Sz8MzR43SsPolGKtJZ/Snw1ZOmAhFWv2QAG2x509
ACZG5B0tCL3Xn9TcF+iW6gva9LwepjpnqlrCjwyFt6Pdk0w7KUc8rnOVhHCraidmo0rgX3MFKfSt
E9vRIuDV+E3vDPdKCdpmN8lHe1Em9yxErRum20+jzQHbbn7Og+B/f2P1wf+eJ3PVDJMOlgmw7S1c
1iJbhW7LOE9qwLCiNDo9jN/Yh7MQ9g01E87ecYcvq2uyOJNDmiKUwF7A19+7FsUoJmJXLOX4d55l
Isz55YbpmTHsJPNq51o8Yg3MD6Qqgd3gO7Abv/S2RXQtRMsGu5+WjrnYn3OjkNklXVH74r3IBVqT
uQ6k5/AFOOhjluJ0vrxVZZS8Nid1fA0M+LB5z0skoiTF8HR94fdMATsCJZfofNNWVCjwFqzUbxdw
m/TSsPIbwFvzYGEmRMgYYkuDiJahgLzeImpRo+4NoGvND/lgViZvJImbFbi7jY7JYekIPqIYbbJq
CaxcdoWJs+hhg61Y5aRsGtdTmQJFKdRrC6tw5sStzXpq4hi4SXZEq3ICUvfhiF2KC1hh3hyFksrn
iUvsxyudIshTbbqc1qgmtK521fUotWFZ/Xne1ipl8GVdfzkN+1WxHU561kiQnAF913hCXvMjz/Ry
BsjXgrMGqQ3FpwOXT7Jt4526kN75jA3ybldSEFXfwBFeLlmyvhO19V6NZLvRkumO4EsBVaf1TJOO
wBEPxrGNLRcP52ZDMxPcxmE+ug0JQ8WIKVnwpSxoUMz1aup5B7I+5cmBeGMJJJ2uvQxSFVWj9wIW
wT2B1qwSMC+zoY0g5UwU1vXtkIbKyVGQUqJl6ESLVyP2rJovacyE8P1n875AWJpySAflXn5vXsA8
wapAfvl/QYOlPW3NBzuOXcr/1q1lwDQnE+jrfC+eKXaRAKKMHuC3uha+p9kbgNjM+hMtnh4jL9+M
m0+O1YnJWVhm7xHVVE6HWxyBHmTx/83wenlyV5zA9nuEiQ3nucrWhvt2xlR2Q88DjdMZO1eZS36x
LQ5QW4CcpwoT6Crurcw/+sOPS3j980d2OD/Wi7CpCn1o0t3tj0GHBJH614mZOxH9ZdiOJvZSWqTe
7dhFxrqw8gc6FS5FJ3Jl0D/c1Siktfaku5/THWLoNXC7jjXeE1ub2NB/IRq00uYuBgUCokGPrsTB
21+yNKTXJ+rgkf2kncTM2UYMElI/lyuCTX2xhUCKEaEG3Y0HrVg0XylOPxhvYdWNd6ey17uJbzer
5F1viKoGM6CHTqa/DXwERgbNXoRzCWi7uoD2zaK+uDChjjex1U7D0nmUG3xjoYca4hZLqNDGWZe0
MLwIp6BEtSvsOZOXZDD3E53f0i3068xZvbEMG8mSRn3EnNtAvjd8dRPBHyesxe3FPd9ZTaTLkiKL
TBuIeAEDiVUJ1okayDO/sbRtF1nUhuYS62HUsVWGrsujKtCmu1iXckVc2Ab7PnRYJfyU/JSMRZxx
ETyKcW23mLkr6grNDEqREa+//nBnMOPqI8o0egFANdYblIXBcNfIeI8BZLmd7hTrgwOWdZA39QkA
pmz3dX+mOrkHxpY9tAJ2ym5ifPyN/jbeOD9blN4K75fIcpw5IU1CNBU07vu7XTGQKur5tyyYIUcz
hZplIqgyFkYBIQkI4130KBVPk9fepOZPLnOjTsPT5iH9Lv6T0rhVONHnAJs3pP0YG2IX7EV5hobQ
Eyi6HjpDSpL8RAcKIlbxXM+tc8me2tKiEkH9usrW1JFgAaY14PTGnWhf9knf9iiMTJLsMg2rmXm7
wzI1SKbw1TmjIYp2vJ+RLU3O9cqlJOx/RVgsiixdxd/knOle9dPmZ5mt0Ml5BJiup0G5i82xhB10
OZxJ+jCspNIIvIpB72T3ui26ux9YRAQ4nDMZO8Ri9PI61/3aZjl4e/vq7fvY/2Vx866jqEPaebwO
yiCdnDzwgyZPkbJDuKCQ5lmFpEyJ2Nkp2sFVyjHqHP9iccEOaJjhXT1+CXNHuUN8OGz8EG92xugB
EBEo+lIGvG8Zph/ljQbtzfB1uZq97TrcnnzKwoCl2Zt5bjJbi7zWLtEknJT0D+zTEM6/06G+ZBrQ
3aP0TEOyMipmYkdBSlcDfSMBSwI4yq3hR8DOVdiSTz9ARkt0VlQEZhiliJQqAVRV15gPfFZ+j2t0
p0mNVq9e0PNjEnM4nl0Vlv8DoWT+hJTG2Tvpa2/K+ejZaPGJuJsju3YajPf0scnvpqJWW+ikJ2yS
+glGg+ZJCT69TBu6+6X8chbSTiNHUHdoS6Ur+GbkMhBzuNKLTUUglwcxoASVUjbffn1B7Owap2DM
47TcBsBe+dkeryV7wWFcHLIYj6oAtAhLaXsLLYDAUb6mURDAaun0QzNLxC7onakgMSJxRs/reQnf
L7UK/bql8qVayAeFZ42niATpGRoH+dKIYXYHcy8jPbjOpHAbrPLQI1SCQUcHe48M2p2IbMf1RMmB
gHMZmlz7hGAn0J1azJAsJ+AYKyXZxZvPIPb7JGKiKPHy35sfEBdMgNAUpv07eRlnRg027J/C9DL3
WMoIwEMYiVZY8DE8mJYBc5DaP9ni3ExRfiI7oJLCmWDJrErL/VpkX3Pu5j0J7qLHVnt9JCtbbPTg
94+DhIxUIEv6ERf5uR+KPwkhrlW75WCrJemEV7EHTU21ip39InI+hLPM88BPz09oo5Clb9zNP1AA
zXCS9+u59YvdZ1HKjWUEaen3qapMjjSM64N1mABh/q+fh5+3LZARA63wfdYaMyZ6E9dPTs9raoWi
z2qN0uJD2VjcCao55oFL7gbWSGmWDqHKZEQqHKrOzIkPfFxBEylveZ6pZiKYMJzWAEjT1GdRNP83
/XUaGAm+B6gXHucGZ7UFz+uL6ZYCTPXNkcY7nf3GmLficp/K063ZLPA7s8sj7O0pknahYwcEXTK3
t5TbCosB8dyFWQo91J1QKZy/5yQBHioJ7lXDPM/eFY9Hq667BKxK0cMOfoHkI95Bymp7rcBxwdPx
wsEsISXpRHMvIUd/6LhoHtvgSbHGqqP5YZ51RCaGDo6Zy8Zcb7fCaz8t6qdewdsJcv0MeUamwVDo
DwC6e48Wnwl3KhyHzDzYlBDdbL+NZ3/IXLQCpVWvGnCs5KwsYQNKQzYku7EyFucbXgJshCXnMyXM
oAhmHeyOZZxUEFCDnItWOMirxkE5/o4eqO5rSNDJe4b7zFkr77tMh6/lW7nK7M5bzn4aXRVeLrn7
kKWQA44tLNz9keMHgxrUHU6lXezxWE8zsvyAQdGJLjimNQqpxg3YxuY+w03m1QebZVPChiGq3HYr
QTdD7NwuV6XwvqgSZGYL8BoPe00Kkfmlqwsqv4F2uj7xVheQqmfHWrtXCTQ1bQHHoXHCH1k4H7GX
W/GzYsVU2ZkLZAwiLtUQWWLTBhRm4dqVlpIm8pOY1bF5tkgdvrjRwjPfdDD+kOhv2nee7pDy54L6
EeOmW7SCXIPVLIQk56D+pQgWecg/hQe5hS1aQ3knit555j7MpOXmaF1KsSZXkoXxtbqionxqd+n4
yh5yVFosl/b1DhqNUoU1X2I84IkuBA+EoC9z154AmEGCyfOa7mh36rv/9VmtiCx0CieBTCObvHzV
PI7GqM3HTkGUWTgY1CKUJo5uGH8NrPLktm5TajsjK5E7h5UfnUKn1fmd3ghWoQGHaL91weXonWeJ
/c0NNty745e3JapLDrY/r+rMMxRp5VvqM7zzDiGPOFp6nm2Rt95LQ0QnwmZ+tAtdo61O5OkKqD6G
R6Ps0mSUqGGj90ZKEeQHP/5wrZUjsSCv25JAa+hhN258DvTWUFAQwFiaQ8uJPZrJKXx/77zX8Axp
HEfzo90/egt9uiPl2JWl0wKo4GMMypUci1vpF80j5YXwqocrVoSlxNOnmCJmV+rIRF9WvovfJXdL
YPBDQlcA3Vz5BOM2OXQyc4AJFUhKYVOIKjVMGIsV/4iHCwQUHgdBVxWYQor5fOWadlnvOdgkPC43
75pec+IMOkkPJwSGeG9t/4HCYvfslorhowIbGXIidxNY/q4whu2kCa/mbLtnyhLOwoI8odcjS9Gp
IWXXDiwXIxXqWgfEjUun2mcdiL1leYFInXzBCi7grJiNp1mZ15TNwaCORtCUBJBqAAeDyknWiyPW
xJrGQm/GIpM4N8+ljU1rKU4kS+sSNrR4xeVAFhgdVS1xhhtAZH5vzbls+VO6Y+KxfAKF2YOAYjOh
2Dn81xNUQAOHbF34l1o5DHwbcczaU+FkLIZpDiKkprzG9Rw5zXP63l+dSWcDt2c9OfGkbkQCFg0A
dHmAtONgHXfVpYvbZHp9ATIF3fg+FtvyM9rPrCiTHb0OeyTFwf4FmYbNpZqt2ukXtuECFdO8/HCD
MgDUEgtJp6Zb2In8r+OBm3rW+0Gh5m7ws+mmZnH47mvIzL+GkGDJBlwMmrGbO0AvVXbBeKODS2Cc
0MlsRT3kW5qF1ANXxjZ59hd6x3RYabGCtwhnUH+CpwfEOCGAHW5LkG64gnrSBCcalIv/kkogiNw1
7eBap5BeECPQkSmGZ6kty0x1E4TvUOTVOpuMx5PCgQ0vcY4MaB3eXBa0mtB5xbKQhEk2WgvMRhIz
nZvc80Rnl9VGPj44T5gUgVS8TKD7v3P7tQIkvkbo/guxt7V2czMc93NTXN3yPJMG4TLWIou2D/40
oyRGk5Q74uuvG+ESAKgJTK5ggeAQiRCLDMelr4WUlSDUADYE/HRJbgAuYoTrlC36inQy1KWPkRA5
A/S/0WW0juTizRJ49Db76nT96EG8vByrKYLRztAVsu4vvuAQx6YOkODF1UXfoJirnhEv52zekCfH
ZbGEaZ1ZZ09W9PwgOWOecIpuCjm91TYKFi9qUde7vDAkfWO6AwduxnH5+qV9vDkX9tXTLyHSVkXz
FvZ/o5WAumY4VJfMVgChNbHTtEuhEQpUz5K/NC17VMLfhOZ51C3H1l5b1ipQFfBHhOFgjcCRtCzB
VXSngpZ1dwo0fsPjATaEffq/nUZb133S5N7sBoWpr28ATMWazxOlXw9KH+onSdLHC86NIj+dmCMx
5MaYX+fjsdpNFgDKfbXlqxSPu/3o3yGY522ZcsTYAUbMxluu6p6ld2qEsq3S5sLHy/f6CpCOizcc
EB92Jz2BGfsIsw/HC3OnvrQ4MT6mJ0GOhf2MHqtAeJ+CMMpXBV5BQNDl3rO0OBpra4CzC/wslNyB
wXCXxVnb9rOa+2jc+172M/fIOq3ce5cey+6NM18S2WaimxfyZ1MW4P9JAJWznIf34GoZEjd/I7gU
ZRcGE2iNCte6beGOGcKZjvwaWv98G3dRmqdAjTf+akso/Q9/F8XU8x8Nvlppb3Ailw316LnEh4OZ
dELX7jf86q7GOJKEfXd/PVXcJUfXGZxc4OeahrRnOBjynD6SuCYLSkeI3o0dLDTGgpZ96hthhdCh
3aQxwvr36fhboh15Q0X2xniQVi02fAcHv+hUPBVmu6i2sZ5szj46E/ycax7wBLExl8b4XN8x2Xr4
YFCoahTU0/t+895ni2imBG1e6hAx3uoN9Rbj272gnlwugyL2olhkZds9oImICQblLKm7UqqalEoE
StBBZz3gqMVTdgv2IaU5MP4PM/p7qDECoI1ve32f4Rr5iHKCoXouetJ+P6okbpz7iC5Q3w/pqHUi
yK+JkMRNS5PX/r7UK2DURkVpVHR2l9VW6PTcMTYa6wmrHLP0Xcox7eLclyiCvVr336edFfuljPYa
mY3JwKS0rRz5FpIX7SBXs8PJp+2haHpfu5DoCc1xHihNXc9qTMbEiqFmRPGgYkYTpE9GxBOSSPD5
Ig1csEgQYHSXeXOU4cUGnSZZw9MN33pYXBBPn/z0zeslKWwup25E3kaxRaOdTe7WY9Y+TEKwoN6u
LB2zhGFHfxXC5EZxHh8zm1+hcxaFPQD2lCWQtQ2MFOKTHc9tkPEySntQJC5ltyOSSZHY2L1P95gO
YsJaiy6rg7ZW2QMJEFal4YbmcRoTMkYDEnltpLwFy+3I7U8flX3dY5dAYNxVXhzc1L8/hNUOmLM/
6xVxPeCHCp3v65MZQdOt+hCeCQqVtoe9NtpKXausWAml8jt0kaLTbUqtTuS+/bHp6jMOBEopSDov
4gNPj3bmRA6qvKcaqbCO3EVwfpGUkR+i6P36nmc4kbCfQUzrSeJrsu2vshMKtuyoHljCZgfBcu3X
c4U7/Kl6D+DFjWg0tp+csIkMPkU9hJu+gcDYdWF6Nh0cbyLcDObwSqRj/Pt/hRlmiIWW67ZEW8LE
2GMsCWuIDzEYExiS6+o2ptqU8jx495nsNeoy7xNXiJjm+S33sx3rHjWZ58JibQ5E+7CXHf2iRP6Q
mwVjt+ki6gnurBH+zntKKIQINq+E3W5l9GvhR62uGvUFT7Ge3Hb9tfcl75iRzRha5duNVmTCBLof
uXbVXMrgNK01YNDp9AZVwcnf16b5uGy7D6D76Ew0vx7XsDi/EVjpgNKMIXXlHtAcw8FmLszu6ieM
F232s3twza0sxtxWpPjSczP9yjM5Er9ZyidoX7E+1VK70zxGYBhrevZRhoPLVprKUDBypjH6vO68
xnKO9LnUJWBgigHOFSB2FBfbj/77Avsidx8cogj59NqZnjSjccaiIEe/F931utc1Iwm3iQtU5cbt
Z7jpAbzNQF3tR0E0qCzrwaA1kJg5/GhvYLn0iygyTmE9rvh6yDYUTIDylt9X4ZnTzhXT50FoEnAm
b14QPStZQGI0eUw/6MgZjKPkmJXIEMbBzsWLuh6+gBokEYZAakwG5BAoivMQGc7OHXcv79oZyOd+
zZhsQBWY7ftQxh1RbMoD0fDjZyg46HKa6f3HpFhytq2Z9M3FgEBdt+5dYB3T93kVL88Z84qOeXJR
YERZ4EY8pzjVR4bC57zLA2Ru6Rren9c0MolAM6jzz36MpzzZTrEnH+9+czfCFsBriQswJhnMkBc6
7q4lqE2m2R62G2KywqJ3DEDUJyGmiw7t2g22XbgW0qhSbbjw495gT7PK9X4y4RsmchVuzDsTKYmU
JAk5pUoadbsCkZ9v/0rclc6snUy2Nhv8S1EIFbKhI7hVC/9L/lxr1MzUMdTk/VKia8k8lK52nTdn
8VsNNAtCcr79TnUJ1CTGQOdtlF2O6no/nUX+uulNxwCkbtsvG9DyNBl8yYbQftSp7YIaRGFDs/nK
w2+a0nhWOPHShFGt7UQQwf21+uXQm0o1OW9BcJpXoaZJCaFx9kKAezSEhf+VjvI0cIvIC1BHFyQo
mV4eF6QyCQChPSuoJGgrKHdmm4PhmWBpk8neqFFNFmruzZWD8VxNVw2rD0J+z1kYC41vtw2oIuY4
ZJfz37XTD6k7JQVCXS+q+n2zEPiak8hEgPd2n1ZE7bGBZmLsQVvoRMxTQBxqz9jVGVelTzAVAUCs
VdcFocYARYEsz7BWiJhDYzo8ABUbNilO1po+DqiGhXnhvaU8tozT+l6KP+6TXDJcfVIhKQ4jMzJK
se36QosOknUsK8gp2NfUb0MtccuEqclaj4fmN7wjgSa0vaRzeYt9v39PeHRvdwXi0DLVRADYYTCo
QGlzFFNaJ1LCHs9zoajovf3iy9j/rX/IiKco/1Jk2Ro0+dMuO1gGLtiB/oLFf11Nj0RPkfFohT1A
aMtTh5WN0p76fg2+NyzHtclassbOmXG8BIUZ9o9UY9YyVH7V6oWsmTodobwMGu6wFYo4pQnJPpOr
a/rWyRu5ojEYC+fjaD7BHzhbDWAAU5EcrwnMgCygi2iLApBOnvYHE8UJX/W32iHMXQ5qFDrLEaiO
LCIaprq7B/tHfpbB1ympzHn5pXb/jsVgrpCbNRp5COnW6KBLIyIUw8TBC8Ojak/KinHw06Tj7jnM
10Voi4EJfkLeSQ+nQAohkeOcTLka4C42KuBQMWzv/m2HgiEEoZPBKOFnZRW7yiJJHBRQDVjDE2cH
Xbn8+3YfB2i1Gp4zmCndK8rwY6cdIG+PaLob2g55I8PLqxN3YiLUKwVv2ZShm3jdBunUFz/00iNT
WgZCWtbHmCak/4ocHj3436/6YtjWPbfVf2Cv8aFZdsUPaB0Gj5G5iu24cnQbKajew1FdzrV5GnvQ
9NCWRus5nfqDvofnDDeFNRfX/L/g70Jnqpq+dq+RxZP3hCDLsYv6EOjvlneRxYsYmxRck5cEx3Y3
fTdYMrgE3k2EwZ0KJSUQ+w5Gxpp3/CIzEaQDAtRjAEebaL7ux0kVcCAmbz1q3nogAQwPY1Pm7Lfd
QIfrI+QAs9hdD/TUP8KNiUM38JgiPDprVpTwFdMOvQbhGbneajIbWro8Ury9VbvrsBfzAFPCEnN5
/qzh1OQXQcQ+ZZItELgczCWDmzQpLdU2suTnCgSrlSbNEcy95sEbEBy7VfKIZpv1uWWbqVPxgtWr
+8djh0bXa0zxyv9Mnyu815CtFU51IqAQq9UQ2SAkuAOXIkg8yAbMp8Cx/A7EWM2Beo55V2Gtkfa7
BECfv843iN8TPTwDDlthBgdKy3JSZXSTVxdSPXO7q34D6rHAxVActUNGftWbiQDK2VqJqO7Yv4q3
p/Zwnytxc0gSK4PlMfHkei4ZE4RxqFkM4N7rD9xFv6vVzcJOuf/ofnDsdAdibI97ETnXhj81TUiS
0YUUyTkfW6LFOly7r0bNGcuK4f9kQXfQPOMR7h3YxPu1SoVrgK4MGU1/xfasrcIoGdUAsjW44vWP
N3Y1N3uR/dTei5a22HvytWkhgg8YOWmgfMmJDXw8Y9IbH1E6gkK6WbwyDnzinn2kgE745ySTOAeF
DLbXVRvbC0riLsCq+vSikV8J3Bi2NvskbAwXyb+qvM/bTtMfmagPLArHLJTgozLWcub3H0Zf/stl
abmd1QnpVpk/p2gaPJAo81htjXh3TeBqFgoNrZNVFEV+zvQBIQhnV7YRjTWipS7GzuG8v0O2YaPm
ckDO7/LJFOTOiG+sKz2npNmyJdfR1ymh3U3gZ6MyMNL/ovMKje7+8all5TyQ/rT4DjGkJdn3tRM1
an42CcymqQaAXwhNTq1Gqg33PrfBCXKTVDg9EFWOMwx2jzFtlFNQYf95C47B8OzdlDygKw+SDjwd
9jZwlyXx35mYL2pg/58ay5PO8JVN6hxM0CMv2VHspW9gRhETdsj8bKlPlm2hwL32wEXCIha+xix8
5fKcB3FJMGAD9zLXAcrDomtvA3Ei1W2aYOvhs4OGwY95Zv55T0phjL4T/Y8v4m80qp5+dWhRNZMp
G822a0X1AOzG5ho7VPJO+kIZYhsQuTLULCZfDlC3KnUcGmoJJCWS1cyRevg60SVT280dZ+lxJ/m8
cvpXrOvL8f/g6xUE4l41pPtrlVB3UJlxtZABU8rGWpMRg9Olv9k3YuOCnWjh1GpI4tD0PNJx7hXo
fc0CfF43EFloHMkQPJy+hxDesxKmtGRxqQBcDeUBzMWMgShsjrTwiPvud2W+TxwhJ2xmN5OSinNN
XAq+tEeJfGMYIZCFz3tMzdMQZXoOA1sa2KudrQmWMjBNGU1oKODKeGn+vFW1htEvN+7maQB6H3PN
HQnVnXbFTGv5yAh2U01ZC8637yIWPW5pFhQIzEUjWilgfoRk3IPsA2mDdYSec7E+ycbCFvcc50rO
MFxSScjKB25JQiOVv+AI0OfsUDURRA2qLMzbA3WNiYwU6SsNT7sUDB64pwZRv1C9VGdPHblnO1WU
wRBseNNBut3Nlt72AeN402tntP8V7N2uY8by2RF0pCaRSE8/zVRWYMEGWLeNFmU5x+LGanMOBABD
KI/HtVxmExkJO6YQN66IVjMET7VQaR4kbff85BNkO6MpQfy2FI1bsy24LUW4o2EtoeiRUEuLU20W
7AoQlOJL8/pMzKinTZ52UbH70r4Jbm2h+xYQoqW04aZ1A0QXpEdEfV3qjwYn1//MfflcYE6v6z+e
Lmm6Axbmsb6//0nE5iuNX+veQNzl/RqZxgi15IRXVT0G5ENdhNFuyGmXL9yc1auH8swrSU7mc0bh
FhW3UEBO0ZjWoY+YPAKlbjgBlUVXUvpOQ+Mxi+GMhKI7MhgrSv8rnc7PeySiKXdv3k3yipl4GkSX
G2f5UgKGobhuC1HS72weGgYP1Ku7z2gK+h9H5iHwgzKVk4eHr3ca/TXis9lOtir46mLp4e0d4rXV
my6Pq3MD4U5Q3O63H4jkjLh15SRXIirt0v2fmBK8kopo7L+IMJ/vWhELQb5WlOSWfIDGmA25w2vH
8KtkxhCjDmcQ9XlBk4OJHUmiyuhbpwWdQi3z70mWEjUrSasfgjEOSq7Hn8wTcldi+0up8cuanb9n
hRleUV237GeJGLD8aOmH4mbrc8sHvmaaOyYR/rugl43yP+oSErRyX55fURVTP34Y8TyNmjAAIou9
dzTLSczAIA//H4QCufZ8pNEFGucbnAgtl0/y6aFLJDPT+IqE3vN+fE+2hP4e1sxRX0lU7MeHQQk+
Af1TrsZIFXA6TEoiPnqm9LWSfV+iqnYQRdy6UvWQC9HFnUY/KpsDuL2tNo4HFftcxeO8vNSxkYVT
qNTv9YSxaFaJvDrkJ6MiQQhuP/+G87BSf5s13cnteJ61NyE7U7qtqe/btjcSh9CukSr2+SsHsnvG
uIU/N9oYSkHPwtCmUubN0EOwVNV7pypO1/vcljW8M05YIL4xvnsE6Tyf4Z5ILv22U4EhFzGRJr4X
A64cfusL7LaIGXkJUj0MOe/JYOH6TeKONpdVtgtG4x2E8wRCG2drqzkN5DVZJsQ2+1Km3OUDzB5Q
QzrFI2wqjvJSakN8HXaTbH3Vg3IANvHan47K0arGRdPBAvtuUxGpeMOBVdCLMSAy23xhZOqMlNqm
OQ7XSRapUGiiLvHnT5xALsCHcm35bQCcdVmMo+iqyaP84+cQ4OIn0Bq/TTbZv3JnH/lxMNtTaHJm
xJargLPe7AO7KASlLC5FzZ0115vsm+/ydm2BK3G2RkBU4BhabM8iPY0VgNMTSUUpCXS0x5ijKhyI
VP+0VqYpwMrCslRRiHr1a1WR1gLneQUS/26uw1fVaWAwt3R4NmFRX0gWDzM7kWu5ULl1OEjI+t+k
S3EU+yac3+03LcEyDpzjle938ZApCyfDSdIMdZ3YtSTT/yq1EdPU9rKmByspXDgRbav2i1aOd6E1
gQAV9BEAF8yMVvDVFaSLBRUd5oVb3IdvIkHA0WRTz+S6DY+RfdAmk7G+mE/q2RrNFTKFFbDKXyPz
CXs5zI7OsTAcCwZkh57y+3Sdt8GgyD3Yvvs1hDgOFjMKGzQAJ0vBxNLN9uKV2/XmPqqjnFsMNrE4
pH+u7n/rh0kcGgblNgWErUmKe45fTq1UVdZKzwzKgy7ut+enMTJ072dvlgf/dBz4ZCeCLvM3ksmz
lWSpBYCJmlYMPccx+teTCRWhIuPUANyRaW2A4Lzkt4yRM3aP40xc9Bnt8/N4RdH4Nn0mPDa9rKxq
OeJm3voxs24PmcxDwyV/SYPyrew56gC+A1pefHmw5bRHjd27Gy6M1wE6v5Wj/mvsM5cJ0s7rn9pS
lW3MuQLAuMloymoyE18os5qH5eUAtEiAyK+wFyT6lzaXzqo5qo6NNkfh7iW49nRV2h2y3a9cWPsG
XnX8haspAMU7HFiUWmjaxvXnLihbd4/A/vJAz/Q3ABktPBbI7/IUFxRKgmQFGq/hyPCVa23FIPHt
MVotF/WJCLmi93FgpvcBGOP6dRltAGdnZ8YoHmpfesn44CQgGzA8jCjg6wRWhmSfGZAee/b1S68Y
Rtrcah4GukoP0noJZl7+/LEk+M+U4XJsvwevQo02rRd+MYyI6twYNOlF4nvKqDS1n7hm70u3dLRh
9IeF4k0jDisp+NONGke8JSlOZFaqtfet8qHJUG23IocUlXZhSasdHzuMNlbZjJk4o3ckRHVwNZD5
UNPJNciJyAJV/3duRkaIwXCGsou06vNwvzsrlzsStQNElbQncnY/EgXnpmaV5d9WB2OeE0pDVXbY
xo1G5VynI0O52TW+1O5qLkNoodbOsK0uSTcd86xgT6UcPshyAkcWRjTy2Iiz6ec1EO1AQ6L1Us9T
z6VLV0vgwfcDgSMhosH5pw+jum/bqICfprqEitbio6OG4p/WbOGU1o3ijxky5XJfYoj4qy5bbPEH
+LRxfMOkoG1PyScCRUYL16JFcLkRzARfKAi9o5+RAXOaLc4mfzl9cHoP79hZ9kcdvkJjv5Vyr3ak
ZPQYknWu7hl8q3TgBsqK1agqUQj8q286Y4Yg3AQBuJBxB90yguGgCaYAY6R4NFQGv/+Plf2e3EFh
cX90iVLEQfN18cJqYO277tPb/hCnOQ/3Jqw6WuYpBEt8tBKfFnBYXbFSusPet5vvO9bcwZjk8jnx
5f3eqQRk1BBhtyacu7DPy+vHDZKwjCgEW53DWtWtw3gGtlmtggajHijmGoeQFjhztlg9TTmrWa3Q
M+UXIbyAXpguLldm9K3hVgWY/IsZFANxallM3D84/QFrkqY0Ku/tG2yo9sAaD1RZCz5CkYaNkuwu
XziOSAiUJlfzYOY/J0sRlgexVzHK4FD9hyiU7fkeueWy/8OzstGqQ9KimKqFibDbLVZsMf9AdS3x
fn8ZkZUbczVRSv9mDKZBBZWvKSmmXNiNDLUR6I6MOQZmcFDGNlLrYCKN+viywFgIL1GdYgLhReXC
s7QZAmZxLfA9BzJ6Ix9hOFuMjrelesH1hjc9go4N95E5VPttu8bQ0H75HZ7FQVLUPCE4aqv1wxEo
N9p9ZhcW3QdOGB5rEzfpBjdZg/pJHrFbCIr1156tv+vTKPkVTmf4jrxZWp8FHBJgnJ2w8NrYjZM0
i2n0aGkfZPxSZ/2nEfT/inCl4Dzqe+J3gepjt6QmaC/qA0ovb43gkSSMrYE44och3TPRtT+5da8f
NfxiAxzUMPK2RqGdw8iKWo5hEXG4umwBFldB0Xfb1uLBFWi8CtD01+7lzr2QYyVVyjUErOjnkquo
AlV7kmZ/1fPfEC+ljA9gr+MAqnp5rqaI10666UvyzgzQ36wFuKvqdg8hzUSZb8RkbfHWTHcu5a5V
XlfhJdgbLmiubITyedtu11T1f05MvJgJxizIkhKbyG+2mtbPVoNL8Db3vFOLTWDUukbxTC4nbuZs
97reeSPFyQqkI02fzkOa6KOVkzzgiul8V2XhMzyZkw4oG+EbpoL1pR97uvPjG5oN7loa102Y4CDT
znLDfh8qPhU6Df6pTATxy4TJ8ilLdhcosAuZGIdN8hlfUtlfZ0gcCYfRcVZZBLlB5nF63TBB8ngo
AE4pbpUu/BfIIISEeSNiBYhZDMh5uNpfZWeN8J1hATN/MKLhutSEAJ0K+sWPVrcpN/FkBsVDk5Xm
WGSzCTNOxg+rsO/8vM0UuGjb0jDmuiAVFZpOJYJuU6D9caUG1Tqf/yo34ryYUaIdoFWxdBaP1UDe
yI3uRSfQlexHypfRY7nhbw9miF1oaOAQjbQ7nyldia95NDIIG473MPgyQZ1zIrbj6etfLKvC8nmF
1cdQkZPyX+4KJB4txnMZursWiPW4P2uFOZom/ZTKkEL/ZbftM0iXQDSCgJMaq/asHINiO6CzwRiW
DZ5nC2ugs++InBwZNQB8qGgFy0lMHGw9ovXu5PyV4n2VbpHuDqb0qAKnIY2EpO1rv60IBghV/bzd
ks5G4hrPKgGjZFxzt8YxC5OMpC4UGdUAu00c2HWdB2mA/NiVDs7OQQRwt5SLtfA9JCqjuOzdsICb
VBa2BnpvdLJ6Wah4GrunDBwSlyIxVM5GwVk1Yyx7M7ZWK2tPH/Vh5by+GtzjlGbTyBWFts99LcmK
hY/JZuNAAS4d2czIoTbKJ05Fi7EzCr7vEM1qgGzPBsZUu+LzkAvNVV32xWVCy8PseixgA2cHrkgR
OkICvt5WBZNkEX7wJa6neYXLWvpSHX3qnelQ+bdVquxAtkQhHCho40w28fTSoVnKoUnjfz6VHn+h
SA9SQq9fHK8oZCMA0M/RFFJEQ0BYTlcRIPuaCcKFPSNdMod7PrOsq4HCIRUVvseaUGt0/jVTBPsC
HWTvgnyp/5hKBL5T0TEbYsbrPACOgtHIvfytKm4RQcR3vpqXsFu0rLtuoaCAuw0cX9bMqslFBBLb
P66/4KbohGtMrrPX1iCuSrWohNKBsrQgKyFc2EyUAhc3TsqPiki1bkMWTUyK3k4ISmYJlHpC1POQ
pC1IB2jZ4oUfy7TDndahTmGgtgcsHU+8Z502E8N0bS4tZt/5NhxdHIZnK0G+EVa9JaQ6Rli4rL+I
/nrR2g4dH2ZmPKC/GX3ge7tejgRUX+qG1lTIsnzdYFYkgG4RWpvodPIUUsiAuu466qWzPDIlF9Cs
qhzvqFPjFqRGAvHb/PAfDmhp6kqhPkuownQT522+mrCeCzeU6aboDBw6ACfP6Pql4KW3fkcnykjZ
qVcUv4p7iwj2u21DFhJqG8BAwnR9Hy0EXZActCaOcqxbwlWesYK1+OWjOeraXMKSSqDk2oOsD0/+
n2UbUbrDGMiWiaiYBOCvbf8byZwEW0wQ6zU+Pk2kMK2YFrbaCu5sZAlpL6e4pMCjLvsuz6o0JCex
zHnQ2+mshFkOM327TGYBqH1xK2PfLlTTM95Eo5dK8MaGGym8sTawEqbu6pbpwn+DzWmqrGsBhZy7
lQTcL89DKbSfv4WtLQ15vsI5UFWWgh/ym52I/IL7FkXTBLHOZr6Hs4He7y/kMLFj4ct41rJfT+jp
dxTgLjsHTGnncXRbYCsqpNilfYEzfvUYNieGIeGCAoq4ErMGmrlv6pSasBz1pPC28k62345RbK0F
/VgRFRE6f8XuIHwWWrEiRV6suKFUbytSV881ZOPQGpwscNcdFis75KWmDFihm++LnhjV/0qiBfZK
djewEhDZun09j8A7M47pYFCp9Xw1I/R+hmz1VFTtw8zyGHBuhUBIPv9SJ0/xdqj4TJ2xvdlv1tZC
VV9A4DTJsxsHGj1vGFG7Hl87UIsc4VerYo3C8GVhPPCYnBxFfKk+P+2lASkRQBFyuxHbmhi72Mmf
5CYRuHf9R+966VVcu5Hzn/NtZMNIgcLGFyApaY8J70IZ428tG0N3iayNO3Jt05RsX6Zh+NlXHWdb
TnUg1M7MszYEONcSjIYz7Zx+Nq6fV7AnBmrF1wRqhIE900kZL/F+c6Sry9cYf25q8fnSmtLbixU/
oSUJJ/vbFqDSeftzmI0g2cTgLRApliut/hpCZGk19h3n57vYV6/jqbp+HinLHO2CAe5UH+VHMDQM
xseaetPeNaOkcyLYwGscOlhKgLVfRLfnLc1aEL4O2RNPqKQ4xl2EAKxknEEtpdkeHDhsA0riK4US
vV6+nyaconVP0AvUh5tyj1Ys0aBNhB5T0Q/FnJ2KtPkliqQM0BCyVf3sk+zL4QXIJ4hEfJZtKHjm
0A/tvtYzVvsPmIMHEvbaYlOHrwv687SIjBO3nS723ucruVxWTTE25hV8tD/nwKvYxbfTQAPG+FRA
aH4FN2Om41afX48xVgsBLSHeLo9JVP5Qc83oZvf64I4RkbtgXnCgK+Eq1oQ5ro//fLl0iSGHrTd6
AMaXXxE97D0x5KYqEtUyhxd60Ue3wKq/plbgNZMlJtkAYMvxyrxNqVWkQGjMBg5Nws0/9IGayUFa
+0honozwYYR9GRz1veligf8IJzACdYYD7DqwwLQZAwTEQfOzzMVlvhm8cY0zh1oA1hSBtz5vU7/C
uElReaMfRuB+NCo0gZPvd2FXu+VZJyPuQcV9G2a/lIkFs71MAEkL2mzktjfgZRdPBwo9GRicBIiw
bnRYhiHGEH15t2omgG0h32S/JyieP1ODi5yxn6t7ITJvUnklrw8h0rBTgr3xu/1RmIFVTiJRKBAh
MtLCFSWWRnKZW9SafetUJR+7+yB36XOdhQkZlNXcH4EQB7o/kKv9tDCsyUaLpY3Uq1RfvKvr+nJ9
gK2io/8c/wkr1O0HvAgxPMJaFOOZvSRXsvviWBMRS7upfjn0eYCWBxgaEZsDU4THKe8zY0plAw9D
evgLmFLCXtrnGMIARPtQFARCgBlCcVEMxrDHTg8yU0ptV9O+nlmsGKFQR5xzMgaf/zuaXERR9Wqx
hd+X91JYi44WaBmP94pwX87p3KsxA+a/E/xpilOvcOYt5kp1sFV3cR541h8z9CXoCQunCm9o7bds
tCE4aSApTMBwHPl7wuIguRuBEj7wU4Gh57mGE4xcpbQrbxGxYpRKW+osEvl6DVxozNtUVIbk7k0L
TABg4b6RZTd1l5cnNJxrxxykOJCkGkEBoH4a6nUFmJbrRQxptgsUcXIkoxkVKs/v84HCJQMBevay
nDHcg8VtTSZ9rvitYz5XbI+62QfzFKsu2DwcfJBBg8YsEKC47J3XWrQsS5gni4VVzD3JV2NDezDM
BV4eLBHW0UykANaKq7xquuVwsYYapqkGsV/w38RpfZ3uKyof4oVUm4m0MsUC4KCCKtvrngIQ1w83
j26OAGc8Xi3xrqyZIF3Ruo2c/QeajCUDfctvb+QwwSOPgrfeN3frwJiaOzQGEp9JFIGj1tyQzenD
4BgK/LEvmR1wtx083vl3QRPN3tbKR7zQeMfvXnZTyx7hmWzoeUfixQl1tmZs1/zZHx6XUCglBQbI
e/MMnzm8ZqkPfNz1+vuVoPDU/3bgbrL9UlNByB0GzyCmuLYPAT2JL5xBARm+gvsPdF5C3NMgeabV
WhhixKMOseGa4XEuCIG2tEpwMTJZ1q6+8KeNbM8kuHmy5TzgTw/M4ip4h118Rk2DVdt3qUI782rz
6bT8SuWMquf2jLYEMaY6pYKxWisLZ8hEmqUGUe/NP/QSA4MNOd2kPnisB+kilUSPPf0hBehFuyHj
HGBX7sMXc50xzWseaPkta2iXMgHcsemod6MMe36iFsGaV+RQdjq+KazHU+wPkgPCNvl2rtvQxv1B
ZrztN088HC3HehpgwM4h0mKUMjf3zH5vllKa+01s05xDEGaPtg5W+6PcJ+N4QVD3cZnnhebtY1w8
2P8b4/CCI9SVc83m4iIe3vHmu7AowtMgFTBwWyVYxoQv5fPI/8WpqnRJxARFor/oM7yHihwdblaK
p4R+EOl5XS0l1GGqf2yBsl5woPPHy3GuaI7wUwRwXDvbxWnNgB9dvSjNoiyNeHUqFS+5CRHGf2yv
6qLOybzKFvTVB3XPHr2VN0EoHOcCKPqA/OAsSowLXogOWfonxQNt2ytGGs+KAqLWq+BUr8c0uGr6
SnmnSkn5D8eDCa/byDPYYknFejJakCyuPpRsrHvtm6vN8jNZMc4zuj+EdX/O1eNExh6/d0vPH3LM
CiN6PG1whuXH1DvHyndRtmydMFlIZVQQ/6NA8enD3RJrCd5NTKBqNNKOqG/O02hnBSNaQD5xUHj5
WkryPBZp7ecws9f0EUmeXhm79Q1tatc+iwi5f4eVMk22YMkkn+5oW9B2kF/0VNrJLEx21ynyHc07
stBpGc520Ti+rxArRGojpCxeXpZXQBDDr8Ye0komHOrBYSClO73459yRqm2p+MSqAWki2QCczImY
yxtcLQ1loDPX2PMepXwUzqoEyBVeQKg4Fs09cJY/qFl2ZzjtjST1WL3fy3QL95hdpUJKBn/ReHBS
ekelC8hsfgDWPaGcTgRT+jKeHAuxmClIlIHzWYnw9ffQ7CvrArKTjUvkz4xR45OHEQHUSSJYHmC1
DR8M+sY3ITqC5oZnsA1zctCCYdSU1/CkH0WtnrYz1QrN7cYWqWs8w4970nQAold0NK9CZM5Jc26s
lplzSi9thYYPbirm2GvGLnLyA6UF314CHY1ORqA7st5EHXpS3AsguzhIje7Z8FlJR5+VLjtu5C+L
+vcnU/vqpbXE0+12mG42DnIT3gxnz6yjhEVsrj+YHZZoXFIjCRrTgWBDAZ7DTJdWWSjB9R8Q6IKv
NuJ+RB9x2Ixa/zvqwTuFH9LyOcYyrUOXWC5HdgJvux8zXs4i0CrRUqNv3nQXj8TIeFEZQrvpGEQT
32cN3FfLETQQwrmc4+4INjM5tsN9xd4P2NPb64/Sn0nr4XEAAV1a/otliMDXVJaUThm5WbEEoi3w
l0eVNSyXVaSZ8KqWypHizvIMKWJycocYd5lbo4Sxd0ai1j/1yWfLL9s4jt7BEoK+B2o9W+A5jWZE
q0keh2tsMqF8w3+iH/epxNllW7jlc1uJnm2lfQU2gbji0A+dci6gtkqlE4AhzOmqjma4GBFVML4k
V9D6vB6jV8FMlSa9a9p1N3w3GoYdUqedxUbHaI8BFaDqi+UKQ3r//nzDpFOWkJKzjzqave2g5lM0
BJIT3dIfYl5AHjFIiWY6g7cQ2zP76h5tyG4pvyZY0XUP4n+GhH4A9jxVu7GlZvauoO0jk7hoY2/E
0jJOQtOHMd3t0zihEnRQbwABRvWaXVWvjNdmJexSseaEAo8EHHT3U+2mTVg2Vg9WWDxsWJQgdyUd
IwvQlR8RkKznjXzqM0wedXrgdOesFr3hIt+H7PE9JoGv/afcTjFpfjApzO/cM/Lj8nTc32lTOwYF
qIv6BIqQAE8SjcK4Q6CTx/bz3AOIiQO7oEPf+3ujIyt78MTYaIhkxTeyb40y+TfhW96QFMeCiIaa
E7K23sv5m2koXLOFUQqXAi82JgLtrkB4ltP6VW3dX2VR0pGbvYFIXMcO5Uh64fPZofFw5uK0kCK2
VtIwvH5oFwa5GV4qKmdoBsJT61oR+JFQOCgD1ikA7I2tnkDlDsKK9MtxVRdC44M9bhVg2SzfstmD
yAp8EMFxACQn9MfX6vRxoPwZql4egtfIEIG5WYtRIr48M0LVQCqN8DWNTCOP7n5abiX6H2a2FUdt
Y0IFaPUfMJsj3+JY1OvlQGmh1p2YPYT3JXks7ENro43dZQcAYy6qcD7pUWrcsTj7XSLp+2cCVC+U
G4cbN183klvcsoxF+awI6G/UqUvJ1C8I6GITryMOweQ2ugRce0wBBnYnjpS54dexXTDtNhFKQTnc
C074ABlJo4tfHBFOGAMN+K/bzL5MGcAE7CPu3WcqfhXbialysJuogQwq2gUONvRze2V+Fo3XKbNH
tONhLPGEglAkeqA9oIOURZAmpdTm2KG6dQJ/xpKaJzFnX8PglPF8Wi9atEjaDOAyh8r7T5HOHgbL
d6Aytq3ueKC4WaDJWrO5/yr1Y+pfQQMrqURX4B1N6XTUxjHOh8eXOM7f4SlsWfykmbD7UBwDLO7F
QqH8oJE5QcoF4ddpn2gGptJKHQRYRroxMoBT/40fSslnM/g0mLsIxyfgqQVtf5704tiTqfS48wyx
wlJD0xbZI79L/l1A/m1NSw5GGuehRtlT9ZvcGZ6KXyRKlxk7xW67cOCtuIOmRJybeoCbGI85gnDa
JXsn4z6OWJaozR/64jPDzbvV9zR4tladb0C+Iz4mlzeWUICpfBWzURQJg8+1fcnYSPTYmvitt6+C
BvkLkX/qjbsHYgodWKuty55OFIUiLN0XzId7ijZ3c43irEEgpcVL3Z3KD9LaqYY8ZGTt72kqyYmU
j8hAO9ELz/hDE7F3on0L7JtiQu1LqpvGqMXpZFxBbz3ire1OTPU8eqBka6lFuGhToWQ2p9ILhIRp
K1FktVV3n1VO+JMlUbmCtlrBDD/BNbDlQlNJOucZkxiSyBbLj8ezx5o/cfkPtPvRyR1yKcediK+3
V4m5iYRIcE05W2z4S3SwKKI83kVljcmRwqzDFTETvZxqs1wPWHvkGm8s8pQy3evAqM4q8oSyy4hD
bSUGqInXoqSDY4PXjwcm7FOl8XqnZT8ikPufR20kFWGE2xj7K6IXLhoL1+9pSfNYjzLe+BGEC/wF
ovsmtqqTCxg8eBxfcwsJABMdX9WbviSF6FFT9NPKs/7aLmNMe/owGZA0dtVGe1HqneIKn/0gJE3N
LrLSHdtpz8nyl+ZRiLF3WxTVBihzsnKHchzONDbAmpqOWhy1H7AKWsYD8KAnfuXqGINqdnAVDJux
2i2txjrSH6MjT0Er7kF7HBD0CZfQ3HLW+rJCTN8WHP6ZQ9JqyJsEjsVnPon+RHkGfdoJyWS4hbvb
tDX/xEuRb4R0JItGdqcTSCeIQea+ulkgj4JQYhCaf9kS+vmcXvoxrFUC820AHQrAXtNPKaV+v1jg
6y3ncy7Ch8am0yVQQKMha3/97sIMKGsLMtn0rlWEcYcfZcblZFIxh56L7lEbDP0ZX5YY1/hcViLt
23CojGBTCKgdWJo5Mn+hVzl9lWHtXv/+rHYsddXFeb0W03BS1bRKhL0bzH8rTnOIyw/ogYmxPPTA
trIlVR5o2yaU4cnFptNmNBjO+8q1iTYsbGeUuXM0skraxu8GZN9rWfInALe1ltfSMJ8GOn60U4rX
cRw+3PQZ5auDWAT3eq45myYCpII3xdxXA+GewrmHuefKO8UsbdEwt5q8zoB9Tb7zXpW05nUsoaOT
S7mbTjgSWuEIE/h8HnbeEp6Elpu/11YYXM2IQND6sJ3CdnfBExXIuryywA6JNiwyMnJzTHPcxUeH
va0oUAXaXPe1XjpGY6BbOTvGOoaGjzfSDI7N5g3KuUiNmXt4aO28vBFCoGwpKqQROKuu+Z3SZ8z+
G3mLN6QI6xqKac1KrthruXcbTOMmSdfOZZRk47VchO8bq0KkMZw5vMjWN+AARw9W+0W43RNuBAyF
4V/BD2VOu1GkNiNeUFQKR1LBzFW+kb3Ejsqa7fKeVbTlj8ZnkKwP4gU2q3uOxw5H4mHtDlVVEDRe
cMyFYu8B5InTnyd3N65KU76trXSjXQvinq3LpUNaSKgn5q6PrPFNYaH8T9rvHqALw07IbDLVJHEp
4+V5ScQ9z6AAO49Hyi0aMvWgvLvXA6xAeUFKlPr3jiFNlmLIUYiFKLTxqRZPGO40w+wNoOHLP2oq
bRuXUx5lml9TIP/QyEOFn/luaWO4Wj0L2QYjHQNmDTBVoucdrcGoxRKq1plbCdWoNgeVjezXtI30
W4vxYiTYcEWf2yY/2iktdRRYUfsnCVtt4Zbut2XODqLpsK0rCbD46JPKwKmjJIiyTYLCu/ACzYpO
ou2UXSrnLOKz+TaoxYF3IX6nRjej2Dv9AssedRU3qxIVKREFF67xiyCA2Vq41iqlNjso77so+F1A
dhqJ1OMberQWF887v8Y6R9gythf0O35sPm5Lp7BJU+/230x4pknCYLHAEGf0aS+JOoFth2SAy7uP
ERCt8VMxuI5NEJycITPmMNjftnH8XiKDuBKjS2NE5hrC4YAXCkqBEyp9OdP5LKXx7J0B9hODf0QZ
lJ0ejHeNKcUPn3+rJPgFaBoZSZpi5JJz6UeC/FnQ2634aZYFbiPd8OwkRKTT81GlXfALkngfTkem
4rQP/z1Si5ABHwSwJ3dhcxHuL0pkQW/lNvXuno/pKS79WJ25f1Hh3v7GO415eawSKFMSfpVRCVg1
IVKvcMAtIevW/7zuTBhT3+hppyPPXJWlKCp7fG7aFWJlO4ujtORtc/8tP2Yj8qh7TqpxefH85izy
b8pJdf4wgZRnuY/4BJkDCkI4/LHkCoQH0cJ4Xc6ujF4jQRQgZK+Qp7WjHjOWs7se+BUYapx86bhQ
7Nm0q7NrcW1bTOP1KuQ9MXWl0zGT9WSej37RpEsGqn6MbLyJwTYG7pdajJfpMYwoQLdq3vnaN/nT
KM2zS9s4fkwrrZwEoqxIuJGgz4IHlQTPlvZv4lMrA3tyjdpO/yMzQObYNoo0fj7DD1xM2razcLvU
fIX4ksDDygCJMWSDzgP4p3fvSZjthlo2VPG1VcgnO8moFWZnKQRvkGjEkw5B+aR8TyLg6MIYLc/z
8xWEPHD7Ngm2b8r2GO/wJzEDenloxM8tQVRZFcCmGY6F1eO/D9+v8LuK/EgGu7AWKFWA3fxDQQ7D
XD45l0aAQL+i8nlB34bDvZGM87RtXGrFYeeUfrW1PfM8w12u3N48ynctoXEQ1p6Wy7O/Yh7fJvrz
yK0AmysmUROjjg43WwhBsHw9RoOYpBzp6aS1wV4Qn8oRp4UwiJyMCozi97dEuDaqVnwFd5GJxKp4
kg+ylY5GfYBfirY+QyUW5ztuXHQP5cf6ptO1GI5dlcb9j6T0aI4GmS1rWaBu0NnuyEK15zs1XzIT
l+z7/xq0vdWUmQ6yv/TyB6LXE0Rq3pUq4TAoD+CWonWH9VMdSkO9jNTT1w2GGbJmdOzq6uwJTvbH
QmnKbJ7ARoSgB14idjJAO1o9V8KH1gXUdyiluMxR0NM2/3iEDKcaJNUetuGchCtbBNRefeVklzTQ
qBjNwtYVuBmzt+C8EYRVHGCMV+0L+nC5m/Hq4qKzTYonF8GQLNs/CjTPn5PGo+wS3rbkpEwfEXfO
fL2WArfEB0qEY9tGa/KwqPMdG4uTryGEW0QdFU4pc/oHaixhkgTzFRQk63Qnhtvm8YarZpmCEXmz
2wL8APR0l1O1C0mHB4wPaJWNddlAYsEdGZsOZWEzbKJ7cTrGJIa4OZzFZ5u7YE2TRoBds3uyUZb6
0RQzZapNtHW2MkJySStTAv5TqbiA1knYoASF/xyJw+xa0NCbzlA+cS8lE40ElKRJrmyyx9zygqDg
YBbySRim1/Luk5d2EQewE9YtGfOBAmI37ab+sqxaN7BGW5oDjwdUcFDegoMOhjOv8g9+8c4DS5su
GPziP0/zqWezqXQUvAmsBy3xe2bKPoTW4zmKBsZqC+GBKCakFnqnI8q44heTfH8ZUmud3+ZjKckx
o+1V2Rgs9HvptJ8Kzx+eJft6wKPd4rIWfcFWsFXBJnP0kD7wJDRNTi9tLnYZDIWc/qnG2cyVhFpy
CGNwUZ3yDXDvLDld/G7CRPZOffES5+UjVv7sm/k761WiD5rwsU9QKih5ytisZG1iABT9zr69SeH5
cbMZnnz3xyRbXSnjHjpMv3VlGRkHiGe/i0vImE8GH7U+4fUFUhaPyX9ZaSxcWUfkJwFG4mCAldS8
cQF8NzSQxabx4PiEBnGH2m5851kvY6sgoz3w9Zd6+DAUk5voagq3R3hzgGO9x8bNEkc4AoR0jS3+
RS1qlsD6L/cfR8ptrzldD67O6NrFI18xzgFy+rbWVxTqv6FCTaXb80oPdStYJjQ24KeTdd3zTSyr
zb0gRZevZnLk5xO//qAo1e6Ie5SEOpRytYRcSu3hKVKGrA6ux2w3vUkq3Fpll6hUugGCpLDwDaHP
8lJhGHhGPIbq0zdPoKKyfzWIIF3kZpifG2JFdCBu1ML+31OUF4tPRly4YRBi/F7kSUqNL9fYV/nG
cXwNzm0axN9Oq5ChivUtL9PdmWqVrVqGYnKekOcjglgkElaxeP6SYAGEXMX0YC0XPGsaq7qjwN/t
I22gAyiu1eDVhHwPbcdgsJd7Xutfvs7bNUz4JFO42nHPwGTgYT4DZAQ5h9/25OAjyOFHcBn579pu
DvuXwnQFKp04sY3akzUbefcUBbNnTI24LlSbnnyxAcqAt3oVjkv9xZmZNoaC8LR/6ZsDsQ6rvSO5
MmYnTu6kM6uuQGvBE9HHfuxRjVa5xjF0SLiaFmLGjohcbqBGI2Zc/jhKWA5zltW5YU/Lbv4HWy96
ElL4Tz2ZW3nT2egaW7PjrzfprAWZjPf+LserSmA0B0kaEszsX5IJ/uVmsfsKItUc9cTjh9Uj0Gs8
MsuFpDgIaM+gIPr7OyPoO1vkvXXb2vhWcXV8zhMbnuM5R93zyqfonoykx4iomA1dBLPe7YTHriiQ
tBtf72dbGh4HHxraPR3WJoIyCgI82SbAIKrQqswIgNskFtUe7gj1oTYzay1nLOGSw/dA7xM2mTal
KpOQJ8Gmdfm1I8sVAE0Yw/b8018tSV5bhgrOZEgHhzs2WMbaWnzFN8OuHAEfjCjOOuGvyMHcW84Y
q3OvcKB4c1S2NXJknLj7vHBoZP/0tVvuvrVFZvuHHG+mmeA7PtRXCe+qN6liN01hL4a/Dq5oCP5V
sg/5eVNnwr8nNiSD+rukpR9CtZPAm1Il330qIE5mKOzpI9ZvjYKN3bfH2YzX/S0Je3bz3Quk8349
OtWkaLjf12AMDhNwccAHDDP2eUJtoYZEjzLFP5YfRHC9eGcBmaldSWXYyXIH5lcqzuet/8aHl9Pz
anv2yANCqeE6A6qMwGI6VSsN+lbimtu9PNuwHNh0WZk2p7x4F2p5AjOMCuuBg2YXOjwYRqEzkZ3u
UEIitCIJ1O5y/R9qKTmgvucbYSnEW0/jCq+ltfYcXjYYYkHP2/+lYsvXLOJK4CTGI8FG+Mti1EsP
Eta9voH2LH8hGzvm8oL7oITdiAmdQ4YB8+LzlPe/Ay+UKPMxsltAxrKlFAggsTpqL16CFmvNMv8W
wk0kFfGPim7BUIijy7O4kvBOe/Jzo9XCnCePv8iGTZwS/+DeVRdWCP5EO4nGdsgW9le5COjuWHVL
WCe3uX9sB5OyPV7rdg0vSc31YG1OLOM9KKBNH07tpvcA/oY0UJZZcoKDcwJfOQbtOniLCuLZUlgr
shxZS1w7I24m5hcURw8cgXxj3RTbSwi/4/NVTyvnlUdEdpkNt114XrZpty4yLsNVw9IsiiNtzHXy
KrThSyiCizQV/1+9CC5zS7PumHhkVhsVJQnVarcOprX2Z8BKvTJTPDBgS+e1C8XMw9j3XC1Xm0zD
y29weUOnrnEoT1fCJfNLqEx0qP4GJc3kRfamvfQ8kixOn3EZN+Zy//faJRT1Spv6Fc9zSHhuLMRs
XtssVz3tRvMgO+Ca4EuKW1XbYTe1KcWRa6RjbzVquF7ps64Sn0KkhMsndRrEjkcZrW7z8YX1T4Uf
3xoz0oCQPRY+m4y1ENZZezU2N+2GsGK2U0h4RCveN5tI5K9hCRAdl6I/uw+Ugs50H4KwyEqzC2Hh
WyT3IWyemrPoz1pfl6s+8QCrVqcE/47J4WjNk3Axemn0TTRxzxkZ/Ua6HGdd8ZdW77sSQXYiYk2a
YNB2+47GkQ03nB7CprdElff5HdfeoZE315EQyAKYxshIAM1gV+INU8jFecPtjJ30nq4m9TGUNFXZ
VNyyIFLRO6JuY0gd5aHgZ22ZesJE+RAhD8f3vuhcjMdxsvSgwHzIjmJbCnws1SPKZRSloo30pgmv
CfOrV9GUu2HCHUl6pSGkVMdFkLYhI8u5Th1tCvMJV+beIvU0b/J4HlT/cJkpa1vPSr7A+5eUUcBs
Iwjyy3tEChzaAKb2lTwoR2gmPdZiYLZBnoxFsDz5vWGHpaPfRMZh4Bn+r3z8ZVO/rck02VQ6/lxo
4hOH/WphDEGh8Sh5AfImmCGaxsBQN8JEvpaL9kYn1w2F8O9U/Yi4fiHTnYG/g2LcEFGt4dYhzdBZ
adeljqLAY2C1ZEe4mdOWk8snWCzuUhSVLcIoHq0n0xSvokse1q6GqhPhArK525dkz/TDBgb6mkiB
tVYaQUErEVC98e7weMX94l+dL70yVAwMAVpEQEe1kuhwF04fY583l9esfb1e/c8Y1QTX5eS6yhfz
ToMTDxGTLD6hVE2CaIT5XY8uGobQDY2rvNRGg8vvaW+kbR9b7RHofWWMmFIJccQ7dDM/c65p5DZa
08ohW3wf8vBY1YHvAOuk98gpnkjLJDMjd4FMeTa6lnkqcLmYagLjhWQmB3jE31rOKjO9N+smn4At
W4rTHeAYfBkuu6hWfoIwxzTnstCANpeLKOqXqVwkSYaj7qpJCbzU0/8adsLCVk7xIjdKUlpCiSgx
E66W56k9x3WhI/l0S2fJb5vD6XY97QpdiFi35tHOLOdoUYSNi0clnFIqgekiGZxwcaAZAewMCIXN
4BG51gOtrRqQJOLxjhG8Z9zodPB4uFqrQXZ0rtjAqOHF/6z35S1qdBe46OxvRxkIqEMhl/RPZ/o+
Hkqg2oHAyFIBeTdN6y9sO/HLXHNmPTblEWFqt5/gYtlJ1gIBsxtqJZanR8G8DpFPGiPcnSq5aA4j
LZ3s6Yd7aMoR+NjmcgCYFIdsmt63A0LX+XAdfbJTCI93F3A8ro2JKFwQYaZaqiL6VKwwLic7NuiY
o7hec2ZgJD9w6GnwLI0DFg8nHxQNJRMldcLqWwafA02qoWkdnM3fAa4qiCX2FmH5BH30VNtKjIiS
bQt41uug2HVJQ5Y3tdWdI6/Cd5hL7RusTm1XB+MsDX4F9aFP2l0uAZzZFggqfoXSKKmbA6pHv1XY
fCt+kWqMp7ayS7AN9kpetbVdagfFHkmN/SaYxaYZviuo5y+WAONA2cIuZwDa2UiS6NYaeEZU25Ig
BYpvWbBpBvbnRhbcY9UPVanvwwJo4v1GB3kQfR7f7V2Y48WOL0s1H1+WCiEcsfV7IUga1QQGe3IT
O10mRiY93QMwNmVc/DYjbHG4pvghudgSBkkNoyCWgWIO2gIdWsiWbC0SlCrQC4l6Pmolkac+AXkw
fEdwApdXidMUfoZlPlhYySjSLmLwFpfeZv8q0Ufqjf7x+15bT/L4mZzBtuUZBhY1OEiFH/6q1VsA
eB5Lx+H4NMZLTBmrUHYi8k9y7M4PnGTEVHp23qsaJzvPfmnMyPyL28eF+54TLXQfWCSJQiHhK0US
uc7f7Cmp9JLNT5pA/y86Ic09359RWPQprOeutV5cYVLwiH/XU/u2FZXNGyXn/2y9MmJGZoRp3+nY
u1t24FMdKWvB5hMAs0x5oPhx95nwpJGeWBFwLV145LgspIa9G0Rfvc64ZAT86AXq8IrpFHm3WkFo
LNC+epPra+p7z7TjnEbRFMTXdDnyiaIdCG1POg988TYoDA7l/NymGUUBgm+vjvRaRI+NryvYAUaD
utp/p0h9gTtJcDenVz55BZhzgLUZ24nrIHkjmEMXQNEOeOeUlCMUlF94FEW1OoKB1Ql4WDUYwPal
2yLolVM4W8kDO8Z+BLJZ+buiXLlGt7O/Y22BOOiqWRnsTsTsGYv5md+Xd1o+Gj0tzNO9cEYkGvYC
YZLaazYshIGkLjSkBNzjjBcX+iAAXzh9d5eIllp+GdcAVl5tFsNERcUJh3lnWV/+mAz8TvWMnkR5
GO1g3s16o1Olu4csGJsumOXoBSAqpn+Le9dsUcA9HEqga5LMATOZUtLojBpxqhcfA0CmYbvFnfDZ
Yr2KYJHxO3StlhuaU4tgK85kKiW4ykjZr4izaxi7kcjkYBXhhpWhMDNYyHoUyHbx3OG7qKkJfQbQ
Dh5EFO1cIrDkxFgfR0oMZvJY0y2JNMA63/HFPOolggDjro5pPPNBLbyHCph75+Y19OAZbVNueGfN
2qbF2Y5yUbjPETqMfnJtj0g9Hm7U7QVAQiCC+/1OB0FXs/RrDjEvJpNUfE5x9qYgnxq+yb8nsfXo
bAHij+Gp+DayOIkJeX9QF26L6pV8+9QmJlr4fBPkwN46won8hCBfe5ODNxMnYRO7yJonaJuAOvhX
HPP12+Y05B04o/L+JbV7zUV36HddqhTWCamaz4eN+hWD1WuGgpzeMxvb64kJjaoE5nBTPQVBKluB
s9b6HbchqQz31JJQvHFgzlSRuN4gqm52qjFeynPY8Mqy702KroIPuvgvLoFf2PQMiDVrgqpHMCkO
hxOQ7F+poQ4cBhprLwR4C7rtesChx28n79l4Jhzs3jWzyfwvAfYIHeHqJLlN81oai1VjhE9CD3HQ
LKuLajMEiuhozJiNDHm/VQiig9N3jyDWkta+ez009f+ObsGRNkJo28UAO0x8yF3MygHiat4uOfqi
Ykn3eKHS28lsZ8hbntbkNAkBoHpW0E1N9I8+KfRXQDsEdB8/IXi13KL31Mox0VLx9OqJbi5UCa0k
6DdyWxiHJVkbEUKwsVlznq7zimHhK5MpolSkINmqyBnjaMI2/Hdr0PsWgCVG6zlhy558XWOvZBkC
ASa6TBvku/PfPAR/dABp84+inbzHNH6RjB6naUoP5xUE0lvEPEy8Q/WTP6w25VjIp4CSNdvcoqLE
O6qdNGpZvCerJ0P8TVAcNyYcczDgAx6htHZ3O0+p23mfJdamh6M+7u9HlXAyLOXmivVqtT+mSaJj
JzLen4EFIUk8JcXOtyI6pB5hhzX1KE2gqJX1Lam6QpIMc7QZZQzXkL24EWRZsrc2Z5/rWnpaezMo
zDeFyYY2BYxt7ScSjRI2HttS5GRl8VAHo9dtVsVxG8HQxs2ugqOZtfNw6JFkqYhN+5yC40qel+QA
HuTfHFtGsVa4SEr63xsWVRzncyL8ut+8EV+2xb1ShnGKJymc1rakUBoZcdQB1WbLTgTbrKBqMuYn
WExTtnKu1bNHVl/AKgKKaUHWQSh43+bHHaoIT+dy36wkPmz7BHAWTsN6gsAHpw24QtpIj8kS/8Ei
62p42lRsb1oeQDpORhGFaGBwGu3wOfrUzBTVyzyJNPMSh2hn1e188jeCVcBX2hp1HqGr7FX95Rc3
0iOb5io9uC9mfE4fpmUs6dZGtV8FV4Mi0O1By4PNsLsmffadN2MDfLgLajKAEpdRqCB1khvNcNjx
uGwYSDgZjtMC4kfI3T9JiMkNa0JJgpPSxxohVsoKSdTdpDP4rUSnZhwVGj2Yf2qt8WUX+DrDnIY0
49xDgjLL9s7NussE1/F31K1YieKoCqmEisJCrHFBTu6LHDtCdtew3174Ie/gE5+jAoXfYEJkU7hf
MpHxi6AQmXvigu197YTSoJBOJDRLMv6F5A+ST30fUolhnGGu4RlTz81dzoZSR9Q/ia7qwHY9g/s6
dVpvYDE1op+/GTETemHIMP2+fT7LdnBLc8T/RAeH41mCr6sqQRsynDKvc4Iw+Xk02WV8entsJrcg
kCIKAX3LOqsTqMw3uknfndKhQtDLxe0K1XcWa/LHRYWVPhFtJ7s/1Nud92ICcIILI6KdaHkDFw5T
y5mk0ibjjS+Dc9SePWsv3Me0tUkeseqfPr6WfeEQgCXZEDXS5LOvzR8svXVgbF0NvpZu+xM95Ndb
RH+Gz83AtxAc1HndXmJLtxNb/6UglfuDTJV+l2R0r88+vA3RF9RAKKxzJiWZCiPXnidE/eoAe6sP
haDWQ+OvKDG6sydNQxAVvYHtnEFO5xbXVWulggS+fizbZ/vDgrTkkG1CokQ1d0Hh3E87g0PgXkkN
vuxvUYVdPic8y1D4Dr6NJD7zACRXfnviXYVHDxdOB6e9S8a38MV4rl2M2SJVdgIHTWxVjPBYgstU
o5gPIx0e5opwHopTnUUN+V79cesBpKWHA8b2hBMe67q+xeG9dzYFIlcQhRwihHbiG0NT7aN8Wxap
Qg+UIewhEvNXmvuCNy8tx8oJZCBnHUnyZXp9NAVtU0jPm+jPxpSuXzhCBQprzunSi2q8oKx3USxy
AkvTUg8hvEt7LNW2NUqHgfBctgk740PJsnVFhmnGNGsrc8VAUlh8P4mOTsJUT6vPcr16xOddMCtr
pAohE9e4gQhA678jBS0K6LmRxLPjcCeyUAGgeDkaHJnI2ADI3jvQw/p2Yw2uO4s0fFS0xVLXeNqC
N2vEN+zInzlLUQ81aiRDtpjsWxLPesgRTyTBDebKxz80ynzPydxb32nowleL7uwyVsYHjYZrcxDE
a76O62WenJVsCuzkGw5t9sn/bE6lY7hvMveYn4GIpgjzfGakbi7QiWaEflaHb50lI1aQ2DtdQfV1
0gN0aaDgHH7xeMckkfFF5nOljB/0qTGqLeAG361g+RsGkSUvukm9aGcOU1DgSQggcnMf+Cr7pqz9
u1o6UC78AwtYvpY4D6ESpjmO5+Z25LI/ONvtormEzlhETTDgnRYjxRH0UsZebZzU4exOf9nKXwQ3
CuQaBuBus1z51FDI8XSdowLqtH83TnHb7OJW+MAr4N7Cxf/7tsBhBHDqNoLNfuoDPKKiFORBpR64
E8x4ppxwSoiPd4eOpjkl5zIN7fYLyWkRrNdcWoKkg+S2ba9Uea9M78wNHyLVdIRtSy6iygvQXvGS
92wFaqgi07rs7dlCqDw7yreoZ2+Y/gFAT7A3WTAywUMWOJg51SvTG89kc9WGtqVKz14r3JOGsQq0
XYECCQDg5IEaRMMFUjUolVw8ho3LZSus+8isKVBZSu8vyzttmkttO/OswAOY+aF60pnXU3OAMgxO
ryUf9+zHMu1d7m7lMoHxhG2cT1CWsLYymxOKm9rPBp1K6KK+BpAZx+tvW581Uu787x28VNDh+aH+
V1jyGCh+qGA9rB2kGBw28M1/Gxe+5rh6BaSJj4J8rrOf+xpA/a1oPWemtZ32m10k/L/Kqga8MklN
bWAxwryhWoHtsQdbQavZt3FFmATkKMLJSXc7KTJLSNk/YgoiR5Ohv8mzKQ80XZc4RPDVWIrxjzL+
BcA4HaKzpow9S24CZ2s3mPoqWdZ2DtJ+lhYymUd9Mrv56Z7yehL+EwZ8kVi4x/+9l3ZAWe/XmBe2
GNfSreW7QXCWvT15Gmn2FNu31M/NcR1tp7ajUaIOxyRrG6S+SZj3TMnkEkpH1M75pn7rvHVShXqy
Ycn3/aLE/ByBZQh9KH1ca76zvWF0z6lNeQ8p1sQl/OOyVpAzEsQkR1kjM2RMBHQYfB8KvcqvgU7n
F66R8hF9bgPMlOITrOVLmKkMnRJqylOx9rZPX9fl4MLKH5Y0IcjwfRCcZJ4PBBEeQHKJNviM49AC
yVZT3RZfXW5mn7IzAZJyzRi5JXgU4uSVktZ4RGVBbD4GRo0MaFW2v4K3Dpsga6DmV7nH0pDWUMKT
EO7Oke/p6xN3QsFtWqQCUE51nK+PPR6Y4388Wur6l6QAJPAe+uZMLaZP3/3Ivj+Q9h9O8DHeITbK
Phv5I7aj+ZitKoXZJRGJbzdi6UDJB1ltGl4a3YL33ALx2JsNO6wydMvz7V9CWBuwh6Y7ZX4bR80b
lAe+HKBZb7i1Q5LoHtQAn92a8+HQc6zuxbXLtu5PCxDxcdWm+R9hMaZDVs+5tMyD0oARxjKDn4BL
qIgywpVjP7wBeuQwN7yKkyiBdtqgaRRQREFgbXxVY1SRkFK2H71Z01W6ReUUHrsGW5+//T1vf6rt
/AxdjTCZCaFZJ/JlYqUdFgIcl+LPNXCnVps6ZNwXpXP2EYJPaV4Y27BF/KQU/XVhXqReHInja0bk
ZQu/gS+3avYqSGKIpcrhYBWSXxH00Y78QXk/6YqKJDuDcHErtDWZD9P86pwhGUeMdw9v0LdR7P6P
gB83Ra2L6J01/JZm7sfuoV3nRrtlqAUeaeURZiw5RVxK+FkStfBMQcIhllMG34uNX3BVxIWhtrwJ
uP23NOUZgGkZ/EYtw8ilBhKH/aDrir/GhHo+99VD/YEbkOmxWXoJ5vevyFWB8fZbvBFEYAC2jckg
GrjOtRR8zN2OYpyB8VC3EScMZ7Sk4biRanY69Oc3fUIrZE/hJuJDF4wMSpYNYz8q4dC8FGDz52Cc
uM7vfCtVrH1TepZhqbNsjVrPJYb/U/ryD/kJEeDBBAjhzDL7TNx6jWVc1Xto29frxBDmfL/aV+Vg
o6DJUDZqWhJvMc4pI8dpyyi9rcClXB581PtIqRmIlW0DstvhkCy/Rp2n5fRscM3Ti/3DLfJSzGRq
GPdKEZpFAjkDjZqjuWscQJ5ntddLr5LNtre98vU/3VJRtHMdZBlFj2dAPI67U7KfrnG/bRWvhe+D
NC4tn6dRJRDwyylAJqT20tBDo3jtIH4tWh7jaV6HnuRwWk9Drcx9QvFc1wPn1XiSE+VPEA5KFJ28
aXA+gw7hdtzlFyN1TvPaFxd55t9eam/n262Ntl+EGxKJAuqjZNOC6YuQjbIKZ3cX2L0FL78pIkx6
dQ8gSVzhvlL1dZimYduixN7YjMCxDtgVNawNqtqNQlnGwX0kfxqh65I0AgdZGhgjDvCNXNrjLfUO
b23zCZJO/nwBPjKvsoV2P6WP+DuRaxeZD171nbBKQB/7LPJOiVmDajkrd+gyBTEkmHOeCMLYlNUr
9i8Ng7y703frYsqmvNU/YPCUc/NUfF6x2Q6qV+rK4SzEMJyVNT8kfVa+pfWY1Bc8baUJosWHPCub
1X9swfCl4bZR+wCEMUOGwLXl19Cs2HQNn8dCrYNjDr3uvK5hdYg06huCgS1qOg//b92wZZS/rLT5
6Q9HiFyBbZmmUttWUqLCYKeVxG54ssseJ6dDOFafZexfMDidZ71KX9As09PRiFem8bj4eB/A4OCA
laIIS9VvaYa+S+n7hRRn+Y1K+OiEROGoLNc4AucqnQXJQxR5rx8uDxu5zOAwd381OUdsgj1eHrVW
Z2cZgtQ/KIOHvQsgaIP2H4FTpN61XvTyzt2zclSNA65YJIiLSBBnHYllycaNyrKWo3bo4wAyDj6v
Tuij+9/D9ZcOH5i5kFGIUmyKVwhrjDg7nB8jitvw+u5cnBGe9pL7YikVQYOCKMKm4A6rdIfbiGic
dA4bZiAvMozSCYj8OEIwluht+v8QXjvDokd5575H6zq3QH3jqYwwueB1SU89qfFWX9cD8tImmv5V
8W25Ajo7+PiJFz1bJoGIXy+cZ4s19wC/6vJWK0q1/Fl+LFparplCi4cyFI65iU/8vdGrOAC7idAk
ise8KdiPMNeOw3Sq2vYV1/FWMo0tvIPFZWO0re8iHJM8GySbRmwb+ih7E5ElPG/iRMjWGzBbxFiZ
MWeF50aV/zyzGPsEC3f0DDEr8FFwlMiZoS29CWfUeIlicKjJTlTvLMgb6liVtQJJv58tOIC3yVzd
M6KKZQ1+XU+gLxVzLF9Dq0jPyP2O/xrOH7xIfDXFd83ptmp+yiA51Js7FliYiq/Uj4u8fg0imOyS
u97qrd3mkyurFK8BONwkSpZBIaRIduJo8VQHQ7IluPZB+Uuq2bwhMy5j5OWY3LWc1jfksmSMahUv
DXb161JWpf1PWmLYTthy8AD7W1IIc5TSLT1/y+0nPOVL8sCPb5tLC8jIpt/KKKpU6LsEH/kzsnxc
WT/Pd5Od0PG//Nu9vNGLzn1O6hrpy3Cb/eit6Pb+emuzWfog7eTrosTGEmTeCNT+MuT7hXYabonW
NeTtige4lFISyS9eoOp6E318cBQKqZEdkGykEnxt8owQHGi+3CeXUON6e802hwXAQrJfPBR1V9aT
GbQ9FN+AgCksYRUjDUzkNGQHRGSl0ZrVmaTxo4T0UNXwfNLJvJN8TNFdrzJia/upUwMc5Rhm7wHn
awRwm1Bqebr/0NbCMKVkG+3fHdTXCgpPC+5oFr6ALtUTn//9cNY87TJySwuKtWjosdPPlShctKlZ
Qkf/6HerPWllqRFiYtvyjlm8A3YtvCMZjfK845kLlu8zE+oztRa8plz3OeU1wteltfH4iTTlKe6l
s9ZGKV9iB2BmTNtFvf6hnc6gFAouaXbnu+W9LulEWLrosdy9oVz8zo45nbxEr+S3/Vze6L5OTVmd
wmd3yydcmdfELnBsv6GOLzC8e7lKS+9BWrpJW2+yTX4nVblSONNeSIhFoGWxPsri2ECXbJgqTfcc
NlEalD3DpgOoVIo7Jtst4JEeTYIGkmFab+IswCbFDQ68KnFrxfn4aIRdx5fZIHthgJhqBys24FLR
otDojFCGB7EUFbkUcaLF0yn8pg91NtGSjtLS1urwc+7mxixnmJ80kivH0EwJFnofZQIeq+suNrHY
poIYvQzbbnOR2LOZl+SyvyOfEd5JPcXp1T2Ju4TZQCCw5mN+YSVwfGWWlCj5ebXuu0vjFhaDtAeK
nas74xTKsogKyzjYnYUsD4/68Mli+LkLEkg8ns84yf+vHcxZ+ZzzFXVD7Uh+XSA3qCDPfwzaITWz
T5yTkvqyjvkrR6RjZQg/mfkKn5L+IZVvdKwTmkGY/PHFQntHdVl+d2WNTGT4lop/27uo1MbsgAbn
apU5FXZGhG23nTMTXc6N4Gz8tI4OgLSIeLiQqwnScVLdfYeNqJtpzA+BtsQ7zJ3Or2Gic6lNmRld
vStJvJ7nLkjUQGMxvve0fl04cIs0LYnumH7amrNNsdo3UdGzVFsURlKsdeve4emmnjm3c0Ubj2F3
sFFsQBQ+alzSdhlH/dwlLryEKczJdLUMa4fafCqW7oeaiV8Tu4iRPd2RW5HbxjUbqTBhjdJHVI0i
mmcTwc2qANYFuR/cPtvLEhopVQgq8hzd3AvtSEBr/+azLIgYDSAwtOmclVtr4z/JBucxdvALKjof
utypn/sON40AFQtkY92J0bKKMvfVcL5C8RDzY7CmYxwWHWi1qR2IcbnlDNmzmll83mGsHuvOfxw2
41Yuv1adY7RtvmIEDAMcEzixGXlzfDidC/M5fKOhroP0A+/4hM615yXXdVGhdMjQbsOdCo/TMJfJ
9XDJWvvsxd3VKStLuJeU6rB8RMaiPvP7hxgnltAt+JZU1kF5SIHS8XKRD0TPsUjhWybIQuKZxB+p
7zufmVFYB00lfDmLlUs2PMhrZ2soU5ZmgecSw2/bgMW/TFD8RqiVMuK1+jugNXNGmLa69g1x+a3w
r0MqFWnZRtEa27fQcDnXO82cFcxOBcrzcBY0sLqF7we+xQEiwO9r053MrXJxM0DjTm4owhchoThY
5fbP0oH+YhoEmSj/HaFAnleeeNJdnh6GLB0Iy/iEDsxf7JsvxvEuIcF1e1TZtaqYCPfTbR23LJIB
W67mGuBF3KKgduS727E9diFV8OQCbzYb3bV8pGefZRdm2giXyjduGz6dLMlJqUXnRiUeEmjFIzJz
x8d3OJ3uwcEcMoMOef/sY4lXk+EEXh20FFxy5NP1U2rZpridSbhZCIwlzJ47dwPmisx4a6EXvntc
My/Z619riyiPQk4pXk96TwDddWSiX5/gocgtOHf53yUv9Pj60FuU/sBKvQDKJS7I3qdVB4aY/LXr
sUBBLllJ8OPp6ibNsF8H9fg6YhkGLIWqSf9sUhVsXQNzvUmBpWpw8TUuuhSCgQEJKAz26lyULihi
DZdeWJX8FCu1H2dDVtZf2HhqBZ2duuCDe388YTz57zrKNGcrKk5yaH5iYWl2bm0vAMCoYCIDUCs6
V6Tl++k01AqZ6/CsKg3hHGAiSTVFsA1p36kSaDoxuGWsXU+zb5f6xyExHLL1DPLnknVR7HhGmgjc
V23DHwT+ocg+W+nCm48v/15ybEOf1rnV/JTLIi7xltaYKUjqRmCGeuPEuPAu/b/sORrwCY4UWxbx
Yk2nuftcBB81d9K19ECJ5YS5mvxlJ7aWxrlvBQoWvLG+W9BU9i1n13nSYCeoCAOeqxB4XkVv+5y3
9wUmjnyzzie53TTPrapTz0JRhf6ovIcppnHo9C/2aFrSNTZVH4M+f8GEf6xwbJBHYpQyx1YgjcVn
whoqJBZgHvn+fqXjoeMYtFF7M+qCzh0gFgycgvXTsojVK47q+tihOB2DMqZOE7MutojXdqTwftoh
hNVQX97csBosRA0ahu8qgyJLLPB2yHCBos4fYd3SOjSysihnTPE+EGNkblSikI2XyllDSdXLId67
qkum/kGdJ8qw9knOFF37BcgIBSavD8fi8ynLfUqbRX3+0M+TPTrhYd7nx5gNUFXIJ7lAsoxWtWmU
+9CBIiCFAghuoR4lJ1heV5gedq36HH+QFhpKQHziIuM0aixRa437Wl4V0reBuivki8Fy9W0HCqqs
w8tIc8rpcoOW7XwiUtNm33eVX7tVoVKtEXJbjeCivYmBmujgnnFUu6OP9yQB1BKkRkp98KG7A4gh
WbiX/wFT+GfFkaKPrWhAvBFguKyz0ULROAZlx/qPWv969SMfeQZa6IvnV1OCDwya+9cLzPOLHrS7
9coS8/Rga0hYq8WulGIKe7ECbfyxz3rwKIoyDGEyAWYdk0C6UMEzqDG02xozAEfHQodBP6nF90/o
W9ZBjT7kfyV2xfUul7QBFkOcUqQiihb7bP8MmafDjcTWGh0ns38+0SfGECQ/K8/4qKSLkjgGlPLd
nr3VFNI1hJVLQXUBS41xk59oDK63A7sLJ1BypMwO4fRlj9tbOvOrFtLRiIhSzv8m7CtinzqJ9STJ
NCAqfvBiw/LYGkfbeZWgQhAvjOvboa1R7E/p/esTtsmrXOvYGnqudVhrcCAy6x4/USAokseXmIeI
4EHj+timADH1siUPCpzNIsJ9o21z5i5xx5lx0j4iHnzXZfsU0BWcjlIM/CBHeA6NeytVFs0ZnFof
uXuHLhGtfnY6wsWY14dQdk+y/rfJzfsHPJnN8WVqHp5YWHi/WTu3BfuSgR6CZttdPe6fW0vJmSCW
Q6atZMvGTdmrnqsw7GVla86pvVcdbKRTI6fnIZy1EiAOYtzRtTvCvvl8iUA/8hvF4P2yltd7Hrgj
EP2gl09xEB6fFktR+Gnnzh0c9oM5skU5+gbpbaPjpHRiXNz5qcSa/myu2tF7nCCsPpKkajPPS8c9
rO+CnXHnTxdMnxwDBLkg4i1W5MosECbzAU67XpkVKNydpybXZ3Xonr+vkglZcSHuJYpZi8Ggl4SI
eaS016cnhxIP3Rg43ZRnZ7Cgc4QeBfJT+aeCuAQK4UNdnwUpblNxOOnMkfnAZYBnvyXFXejTf6+j
mbQBzUm0MmGqufUpXZx8H1Ayl319bm9xBlQXr2zhpoJSr/4DrNXUcDtYhYRDsL657Uf4OcctAj7I
iZJMWkE6Llau1tYLbKMpwKHLZ9MaOQ6ISDVi8y7G2EhCQRqt8+oBKDzfD4YlYh1XJRiMTtb4RxD8
ibirO/1rfsCuzFnfapeJdp+gFUStNUTTh7x/7cK6icNK5Ey+MkLs+SGGN4RIYTvSfQcFP9XSH7R0
+yoJRbZS9lEU/FL4Rr4dxj4clKkn6KXTf7kjMblh+SrFNxPve6BU3/DRbxkhOoYwh5++yg8XcGd7
a9VgN8No8xCtomPsN5EDx3ziZWch0wDmOP8ZuHrhktCS/XIoRE0zN9Ukc0V5rg2l496lFweyPWAU
wCg7NFfltBsDbFeivZL78G/Bjd+1QKzp3NBPGIGE03PQMBcgpwiU/SjpHw/9D0xldf4B7nG4L8Vc
G+ZQ9Ds/apuaoA6CUswIfsOYG4BLJBxQuvb3jlISdImUj6EQ9E8Ideg9W0o4WxSuBw9FdEjHLZ7g
eoARHAMeEqJkxXmbrUL6xzEnNyKZ6tj3YKiLSRatYGXMljlWj52VqvE9IytVK0Zlt8WpgIYsRuj2
xRafaSON6SKPHxf70Izu4J1JVcTNCyECy7teZIaaiLH7ridenPHfGOm5ODiwr9figakw5YA0G4dI
DLPksnJD5n4NW+am96u7RqO7gYCsEYdgc38Ghz+blOYJkA17640Wo5Xkme0wM24g2fzFC9499oDP
j5oLUuzxB9UeQg8FUPCjVa/gqj9nKGbjZku+P1Oe+UmeVB0RsDkQhMAK0nSBnf60BB0c/2vLHkrl
Zs6cdYjkdxEBEqOnf8N4QGQcHuawSKb4HQPRs0Tq621Fa6VU1nSjbSJydYQ4cFlIye7KcBWBMJwI
wDDrvrexVNTxKE5eSxEHBpNZ8Gyd+K2PtmOkEItELBshMVMMGxZYIfNkNedrqIjoV/n/N5mCrBXu
NfkmKGNlC1XdjHUQJbLNxZ43ilMXG1CV/LQTNGsHkpPgAT9iYR8IUDGV7BklYwpeX5T4zbnZaXvu
FY6eXkxRouZOTGoMWiF+sW/MfDEL/qvKFvrurmpRhPWSjunyUglWsW+HhhjKIcsleehS+SVTx6sB
76cJhCLQlMeicCpNEZTm+vTRc1Bi1t/3UEBV0rUbYEnQey5tZg7oE946jA91+w9xie7T0FvWcJB9
zSGvuV8dQOq+zh7pSzOH8Ziua/vc8IDg+jduvmhHvVq3BU82wSaowuotQuN7wbKhEjddxXcaAT1c
Fv7ifDTHLOfBMZALSJmz2UXrrERspi6CBA1kNVnG6/LQjBEHS0jYzxubTDusu/1MuvBiZEXCmtnc
nXe9+b+LKUOdDjH0ilPYnB8HK+fATz/NrL3H5pwnzaQqUrcw/I45c7yCoOtAJJPLNqAN+Cfx27Gt
iERxR9AlLjGUDGe3ztmcuV/UmNmeH99sLPfKE9G+KAqgVAQ2GXdOca2pALAnt5dZrAORiaC/u6nS
E/TJtCe7hsXc70qIxWKZU4mfnW3NBQ8D5D0NQMsZ6Gef1KoFRA0uPCoRonZGwNXbe6RreE5+65t7
R4f446xQH7yDfZUp6f5kfR0mw6JdqHqC8/ggegpULMS/6iTW9h4B0ZgFgDbk9By2jwV10xp/bki8
DLsW0c4d+/MU32m3zmIJjmAk6NrLmuSB716ZdWmUi6cnh4J1JQadAHtNfSE0Vqrmg8yK7kYMiScf
ZtRrILENsds8jk8/0a1KY5sl0ANJPoZ4GPwun93QzzdeeGhBTdYkjnAuUmBr6jixwysyO/qB5Wcb
TZ/KLmQvpauEX+KKzS4Y35IEQBqdN5I5N19wvL39kbeXpyBXfIa5YeUEkbIh/aJMObkjyxLmKCHV
sSrNmost1/N0e5+TtmDVddgfoTNWwds4Mg0Ksv3nLG3i4NvtMBk2ejyxLvpQotnbdXzPgKwDZ2BC
DRA3l9zAje+Bnvq6mh2xZWZ0V6kkLUlhISewHlT9ZiU/qsjWkl2+PagbGp2Iw/GqGo9k4wjkiK3b
60m8jgFDViaDhL8ZkJYRNBXuVaqIdZCEFM6Ov7gYkuMSZqvJUHnean2m7AUxzb2VMSeI4npi4yf4
frEcsQdmZDpfIZjTS6s9OBf63JvG9p5roZXlVBDf6YCzabYehRmo/BkkW/yLaQ1krYv5ojn/JN+D
SXCciLQrfFVXxjBgcbtcRpzt0lnUAugSk2dQ53WuCWIqMk8VoKVkMwqDbiAAIvUIUx2G3RA10TXq
Twobwey5mssVsWX8xH4uD8XHJByMciY+Tmv325Q7nDtP9LFsFyalSMIorooCcjK44ujoJ3cP2vsg
euXP4YsJqso69wpUCGA2x2d2UE55z2z0RbDy6heZlK4AnTWKQ3Kt45FzPn6Qr5hWXSMmRBYppYRd
zH3m4PxelqHZtWvFDmyMV3kqznHGj6G/j9gGygeV1iifIw9SJjNJ+xpaQTAVSiVSEVonJWHGZv2b
syaDQxOUm7gHY/tP/fqUWejPtk+cDA3DWhO+2IWOcNPOsPOaKvkshyNHa4+P/NMODMxpvxf7wboG
3IY6hwgyfdSn6vkZVsXJp0QBSW8H8BULUmCOKacGhOuFyw3ZQsXJ6wbxAktsJGupJfN4DytoQxGQ
IJ7MNJIy5rY1qkynRa5osEC4hk+x3mLeuJyNjcvHvltnUGQi35aG/9+JmCcf7Vwgv6zVdP6XeUBG
HpT9JzAYteJHrLDGB4NSThD0Zwti7UTvHlcXnfGVNtc4NtPcEW39yms5+WBCHZxyMtAKsoPoS+Sm
Y0kk23e7EpZ386J6k1QvvFxx+ndrCZYN4YripS8+3e8uGuPo/stAWmACLOTLBLAsET3CjJkcRe7/
Vx+rIMJbsV8DJFz7RwG1MBE3joWMLFcC5C6iF8uKh+/UBZLy/VUj/Xp4Ve8L6fIo87GlPVBXwM7w
Pqt9xDSgx3yPPDS1Hrn5ONurm+Y3xTqrCSo+yFnIiJs+0Oh02dpSPR4/p3mXa/9FCaGQ3+JyKOGm
916FcrKg0JVJRqDD1opvuU+fIWCD5tZ8Pzo95el8XaPRlBbY0hYlfw5RpCrfY4Ym9wBHVJdp2gas
/nsQZxrg0E9vPe5ijo2Lg/dG9ceP25VW9rvol7LPYbRxkFSK1oE/S6cOIxNcKIeejmQgOAC75XFI
hw6TdxWnbJas5p8v4qzSokItPmBKyl/wT1EQz4SGNxJsL2WZNtzkYp0fr16J3KlAycjb/p2nR+Rv
NqE5q3arhH065MRHI9pOmtv42vpSQxtnjMJhX3C3urCcyM+KTbARD3V9gns7oq0T9oDm6yASxXDE
WLYmbSKnru/Auf8vF436S9ialZ5sulfRC3Gll2+7FgAw+kFqD1LPH6HJzmUDR2jKBo6lctOtdP0H
nwAjuWPQIQAMKvREtBhvjf3fJwNw5i2fzWpQlryi6hm5k3ZD1KjZiczxzG5B1irueWQEFEwdziaN
omN12hD6sWhkLHfk4eZgBQQus6BsGHYUf2E3kBd5SKc8pZNwsveS9wKN7AzmkqPMzdGoYf6MlcXS
xgI7Jq51oO2CDjmjKIaT1etd2056i/gW41pDousOehPB81MustOYxKC3TH72waq5YwsXxGajQOId
wr+9t9WQQXUDDYf1ZQD3ecDYgs6oHwTpdcFAHsq2cM2SRGPt+eXwclWoVolS3YnJegCGYLY4CeV9
Wlwms1nRxpmYuGktUOfjEvke6G5ecuFEejYZ3oMIgUuP293p4F3coR/AbwVhvcn212kd9E2SaTM7
n4u1fh70GWn1blBAWB5ARAlCHihkUk0f7RjVzTdrCGpHTrueLgN/gN5DDUlgVUrJa11aLjEUeeiA
guw3hHAjIlw8KlDOagmk0jMJ+D637esUzrl1R2XaFHvj0jVIrQxlzH1UTlJyInGtfmmluUZxspe/
I2yZXwlYn8kyxMpiggB97FldZ+rRsIw2GLDyBgdepZ7QNLA/tAMQSxnho/5XWwb2Y92owl5EpgST
4DVAhoKQ8kaNbLE67FiRjCn8x+Zfmxepz6jWNRZi2mWjD+ABiy6lwcO+1SEiZaCpyxYGe0T4BjgK
kLYbha7WHzluhzouwYT9MxrCm5hSsmVpJwkQ1/zx2uYHXlUBo6+m3JNWQsm/3ZnC0lR6EggOmMT6
Y/lO+7+oikMSWeDHn8+1Ad/xSFkyO52uujWzECW9oD7wogPtYaVYaVcERX0w+yAygeuWezcQ09R+
pLA4XyITA80slZRLHA6R8kRQpFiubmSpMizxwlbXIEXP5y14fHMoTgTc8fguhLZhiwNPbfKSbgE4
igXbc795GyzWSzroxScJ9v7cTE+qpMJO9QrQH39kAe2HZB4OYKN4Xy8SiwN5O3RX4W2DpKtX9hHU
KhF4o1KzmueTbGjTE1Fy+Ns+BtLX1YW+88+VQASARB3uGdCdI/vwOs83iiZKhtjpPiFvF6K9qOie
c/chLIky7Z0CKefafaQtweG4KIh1xPHF6IlNUH6rgBhPO7BMcrf6YTW7dXndZZLs3ieGX9pBuLcl
A47hQlTDO9TTRmgD0/NRAatAus5lc9jOYf4gH5Il/oLdgKReDWEoYxHxkWuG91f/yRd/Nvsj/uNj
RSjj2eJNbQ3TnFIjANT01JfEwgNbfxJGr+YnWq0OOPCL316qXZo/urly5gE8ajYw5vVP/uVkKPsZ
am7twXiXr64mnCFGNKSMiXCcbZ9EW6f9qLytWPIkvwO3J6QpKdZSCTkaIPQOBNYqlWjfGIpQV3pS
ZXe9lKq25jHUXRjQ4maT2s50PTRlm4M/ducuCgASXnvmttd+4DqeSjafSS6K+ACtlrWOVnTRdckE
A3yHPeb6PL66BnxPyapWscC2GkcX4x+w4xpTKMrIcyQumh9EFcp6XkhuCspiAkPa3VLG61P6iIuR
g6NysNZSvyhpdEFBRkCm1Yi4r1192+xmTyrIxM6kejWdymLpCJ+8S3Mm9BqpZwIsRCzp8+9m31dU
V1ZG9vMUOmMfi77vtRjzADrCiv0yxZeDVt98Kxht0p/83qoQnwPJY2M1bRLVT73bEUJULWB375Si
XNdxQA0/cW6fswieDadr1mKip8uf7T5/4HSKMd5ryVNGe+NPIQm073vz8tgp/oR6g7CTqp3iPBd/
x6hP05L31mG0X0buw55m/MlDkIwc3caNZMjCloqhN4FfYumnBOBmY5ign2aRR80Lr3E7RPYszFwb
Qia2bJ72QaxXZRTJQp6AzKiBVTf7furR2VeERNdwWPwd1fxWUAChZ5FYNUhHfwhP6ENtEu+WmE5L
WJuK3qlzDtrWm07yWgMJNmCJCCyc2MFkNR6z6sbKgdIQ6lbD0CEaSRJYU2uDd/S1bWRaQ6tJfTQK
He3G1TVZnL2D5FbScHK81W7F1lWNR9tIHqsa71q8zBkUPK+m3rgUcPambxHkeMBsszn5UfFlNkwR
xxLxx/TLcyL2YNrHhTJa3eoxIgMlpzUVcMbnnyIp7wF0QQ7alupySWwhDIN+cVKEY+cZw1wyCUKe
JgJmeSHvYYA/bczeJT02eNniCa9byqBm0dIEvFxv44+4qfGYiYMvVabxa2x9w+rmJdMRszrVya93
HRH7Z7EeWlxJ9GO+YMPSfNifs85CV2zYi16ZCJKbjsG1pksPfSt+kwr5YS4MUe2+MgtSZv2zm+OR
5jbKzdLt7bmSaithyFGM01B1rZqMTxqO/6RbUYlnAHYUhtSXn/lvmjovSnnufInGB7pghMIq+mBQ
knAqBUXTp34v8tAo6IodhsJ3YkS6lVHPr5IQfAYqL5Q5EIJk6Cud6TpMG7O/TuvgyBZoDb3wIjkD
zYznffrU7vG2QzGIEFT4zzonj3zGK7HVFAqosVvUvQowNxLXGF9ACeqyxuuwyaxfVWTPBUaK4qXY
fICUKI/bvFePsTCQFEj0sorMTv1pblgci1gEvLOfEeYbL3oRCF+1kqneG1ZUTnBVyfjozbHwmu0+
ok9JG3s6UPrVKxXZgd+QwJQY5n6MtVtX1Z2ynhyDbdAWFCOcAoReBCsGLoiScX0y9KkxYBVJWPVi
IssNTha6f34meJkxMu/5xaBcQ9I/Yy0A2hLXRqEUqF3RJv+K69asBSOZQ6LwHgIwChkpwqIVb2I6
36kOu+bNWDP732HtjV69UAmS58EFOSyHKmOzB7qTh9NDfeXvCFCdpkpXL7EDIqIHSqj9R6TzL46G
b0wm3l5F2K7X/lGRBIu7DDlY0SNvqDVQCjKSJc/jlNwIx0//bv+DroL2+KRacbxqKMvZjh6Xny0W
+vylq1Xlb1umn3TtA81WXesPp+iYxu+rP31fghbySF8Kh3G5KmPz+/SQqTXyuKyRU/nnzwh+9sLw
00HmMVR1AgTzLZdCVw3Bals4oYmb32QCrzcUVpin7UJFo490qfPoRwVoYMGrq0VOCyLbEURQbCdD
nv/ADI8ATCyYNDTPEqe2qC+AgKwGqCoN7iIj85U5R0ZoEZHJexlLn+StUzg+DC/EOR1j+HlcaZPS
qycv5BImdelbRW0rML+J2fwXc6IheG8tibiZwwqkrJ3ZqXKD8Cm5wFVU+KC0ZNJsINYkU1mC0PV+
av95kHMAXGmJdcITr/6CD+7+P4s4M5EuATxdt/SqxT2s/ZoJ6YQRCAjUXqSexkKbHlzupDCh48kk
tJe6M6T0xThFs6S3Jjz8jcXjz9a3Clrt3B/HpYQOJt+EgN0L2LQHwCC84ROV1ROz1ypGaMxXzkCb
zwhIcROLTyjwYj3Gg9bql/iTWgobNE2e227b9NeGI2+XYiCd7JOHfcRym7H86bdOt+joBcqKxSmF
g41w9Ma+cTWhJjYZCISczV0R0ncIccSobgrN3rXMSE6GkkAYgH6neb5+4ELI8AUCbvTXLufcInpe
1RJRYF2q5hyFl/rWxEZ/SSVh/4281elOluF9m2pftC7yP7ZEhcJmXB3HTRbU7HuW2KXoW7APnVvh
d9CfH0Rj+BjwE1ChaE5dN75FRYhpzmTRdanxOx8Ja72XzC9schwAh0aKmIJ8Fq72P6hVBdlS2V9q
Ah3TDPUeioESVAnCJjsRLfEryXNxW/p6piN3THroaAOAo8HCIWRIni0eYjLhT3ejZ5hsUYLEsgc2
MhLWr3EpNfLvt6B7SotaMJiBAEejKEMOndByn8GLO0dOllFQfDn1kyL5Ya6hG2W7EHvTxn/6Vzps
0ygRpMkaNywj0ZSG/L3a7rAq63uqB/RYvHsIejsvXQoc0EAay/pwGOeYI9k9+lh186yNoYx08czO
BRQDxWmI+Va1oRf21zA06r9szFDS/xf/JfeMyTXMhl73jxLZtVPDSbKdtY1FItC2sSszLr7lDypu
zKJEKF2lB71V28BfFwZnAz06hcGXEfmm4LAonF8Nrp54wBYY8YuErDUmn13E/Op9nEuLB3EGGD9Z
aWQ3YsQxLCyJqPsZhWuiOeUxUJPcs1YORWguomCCm7A1KIrbd9qoFUevl8gWvs9EQzQ2RDl18CU9
cNtDXyd3ja9EzWG1sQDrDNP4Kt6U5mUjv3uCGncUeja4sQIBCI4+O6yqFtOfKcot9YYK/e9H/QPm
ezfyai3NsqXUA+27sWep6V6XcLdkTkV88ItFKoQCd7stkGZUi28gxXUXgttBJYZ8N00gt5AnYBpg
2XKAQLsRPA12XhjX0nwGQ2Um+XiYYnZZ7ZRyYuvABXQgykYSihoNKFv7RIW/97E3VnanTQWAetAo
P+1kjfzJaDmUkkr2DdSrHuGvEqjN2kIJ3tyujBQ1QGu2AxV1hOVwTnyK4Y6ymCcGK7oa+mCVAPgC
au7KdGQWenhsg+LK7x04moAcRzYgHpl5bJtMygabJraWbH4H9il6uQjklso3dIImF2S6mz8oT4c0
BoOr2qpOyYDervTVft2wRjSePvsEL3mMn3Gu3Ya5J/wUUxlOxH0d77vnf/IA1J8640LenVmX50pA
S13oQQWNXsyh1GGQ0x6VP7CHzuhr709PjovGnsp0HGeTNtkIPxWTK1voY/E0fPzuaxuRA6g7vK/a
HTE18DxOgPjxJqk9JhD9470mvm3JDwxzv5LhRPQ6Zb6QA3vcWQuGHgC1kBym0nlq03c/kq7teKwe
yB35Ti5b22/CmgO5EaJwLHcGJhJUrDF4GoPVYqJs0y3OG+6Ipou1idGn6Re9lcYj+JMzDDaLJnFE
uAS9k2Q2T1ssFxGXo9DZU1qPUzE+YYgnJdr/pXPU6fPyz9sO+Oqrs0zJZNCmKev4yyKI/tNyeC7A
PxyDgjB8fdTgMHbcsg37EELQyBdOU1tiBuO0NpTySgtaM+kLGXAiwAouuZTMbFbEKAVEjX4CjQIM
6jZNpJg6zFDP4O012Ml+0XfYaWiaknVhakEpMKpk3AWQjD/WeXN8SL4iuDrMjA4R02ZNDoqDCexN
Wx3kszbl7Z17kMFoMPagmmwyX3dwmX2hAz/NEn5PsS3QJu56uYp2RnkIysXFBigi+J15Ow7NKVqA
TNlfEILF+g+5+ldtBEfubItLifp4Tx3CN4d/Fm+yl1kZaAoAYzxwkcn0+4Xr3TwK/Gs3tLj+ZHGz
tRy2RzKKZVcCYcTN92+S7k9PTa0izj9Hwhv987faEV/C0cb8d2fhrcaCOXOY3L5rzk9ppGvaUDAH
xNOjWEoPhlFr2pWOPCGjUdOAuXw+saXn4Kqf4kpoaWhoFgoC0Rz1lsmRNTqLWEGravLYgZYtO1KH
hh0RyxHuJS85RIkiJaLZgzgF8Qxq3eqR3B9YMfrKZQrtgVFqb8+CMrpaUnA9yqgvDUub/sp/ppi5
TVx2DbBDAtohicafJnHPwjepUVst8tpxnTjui39KED0ynoGRI+YRhV+0gOxVxVeWOkrdSpM/XWcG
Q9MqnGGLXXoEO7gcZxeG2GFfkvclauzemTZlemMmgORlWcUSpnXP9ovRbp97+8gs61JXGnjiVRVT
4UYffViBbqv1xHqY8m6fHVaSGAkrfzQvZbr2wz45lKoGZx3wOqkgyzcQTNppCJt3xImtu3qlNQnr
LznexC5r1KWpzGmZv790XVaCTsulWPFd5z5PTwBZ1h0yirc4Jb5pOXRG8lQo0a6s8RVdhGm330nn
CoyX+Z0eJOu4PyT8Tz7UquRw19gCN+SflachRsRQCqz+gRV7aUz6lzaR6QlI9gftbu9n1Gg0Llaj
dTOONMAJxilV1CzsBpygfDyxYlEhmsi9unBLL4AIaoAPB/MrX1zp0l5+h8IhA5rgFDn3s/evVMDV
pYMZji0HsMydhGuNa3o/4qf/2vKcMFypMAbrnT8E9AkuH26ByZKXazS6nY3JFSb/4Zao8eL5Zq0E
4KXzrvtb8506IhRwXoG6c9fCaX/VBYxc8Nl55xL7y3Ou16r5SYvNKIAT/LoMsg6MQBmgWRfZnONQ
uk2TRtUS8OQ97BMqaMniN/xm+p/YKixz1zXO70cXWPOK/2njS4Il/MxzgBCWQhP9tSRgy2vnAGfs
V+kRV0SE3Mk3KFWRJ8m2vnNxF/K7ci973UwAqsckbBlD31E0mOEkB4ESC67bARhcYpAcIeQ9pNDD
dsD05E0quNSH5PXcl6segMywkueQgtKZxW/syZI8ZikRC7ufyoVwmmzZ23WsRCgMiXtlwvsdU4nU
bMiWU88eRBf7Wm1PCAk87MFg/dZQdkK2O3sUQr+5Tcr51H1iOrvr6R+pswdFqRGAJR3Ik8988iVN
DAbt9lLge9RqSxch16EiAQfFZ4oRpgYpmFvRsExlkNjRc4nR4kAl5x2hnAabi//ioJYjQl0MiTIL
r+TBfLfn2xp4TkEuGVOz9wEgd0Pk4QXElSaFAkvhkXeI3ON45TFe9J5PmBOKn2gh/dBBf+zB+5iV
9COnWdYojRsBONCv9BH/ahc36m2MTfx0+npKnofgTORAXmp0QC0TxVLfL3v9eAwmSd+YiXyrJ8Ar
/nJmcqNbORdPPHt20c/Rmf+Yt70HhZlqHioGSqVHJotX1gfz+Yx1tLkb3JHQ6BRhB3tTTueQYpRw
wuCkPnbbp8Hiav/iZmfsD047cp1pdvbfPK8eBXeda/vOKMHvoKZtrghIf9NxxliwLB6MjwLKC56Z
i4rQZxIzCwYwYC/Rzb2139n+mdyq+e1+axOki1b81DRwvz4qDAG8yDPH/rYkFpwlCm7RSkcJnqP4
dIDielBxDTFPTrW4pEreqlTqgQx5Nq+ONkestkCvigT6v1f7c30HvcKfio5hqENe9wkW5T0gM20/
tE7+gz7EimeEfRQrcCdFS0UFUCq+TF9GpeFlm4Y3Raw7VxpAc+luoYnxEgSYPiQCP4p6QtaX60jz
bHxemdU4EQTKhCvUfcqZb1j8LT3aGPQMNhGvDQhbLhnm7f/ri75JB8j7K/IaQyIvmMrOV4O1b0Hd
f3kGCCHNPK6YY72lb8hpG528RSSyjsMHs5LbZXHArYRgcT+nuQxq76GvPc+CQxDInD2maTvuz0fW
h53jgPXsgmHNOD56Bff9ToK4AV9vmenNilj5V6KSSKCtTqd95JwXagXeKlLMVB5OdxzxPtOoBIsf
Ua7oxICuiPwYmUQGm3pds0qE9Aq9qIxQebprTMCZHM+yhkWU9YNc4O52Q1EEhLKr7UxeJaUzkhoH
DBVpx8zjMYn3aTQOGL7A1qQQWFUswZmc5ilx5kB/ZnkYHeeORip/eThe1ANhBTXoS/wLDAdCJgvb
0LNDi3zcRtjIwvtBLDc+Z/zxUty3sWLAXofvZuUw/HRjXX5ZLO4gNhrJkg66U0moFKj8aedfgMu2
COC+vublSbpQMtNPKe0HtnK/VVOIzkAxX+w1KTe1AtX0KxWbqdoDgGx+hZIZ1TVoGQMtqyAc7x6u
vktd/1Sont+KKPnHqLUyJv/xo7D8wI6IRYu6VVzdUCDk8Z4pJ3ONV8lCKhPEf4phIoZSoZ4+/PI4
2G2wXDZ32rLZbImCbztFynjInLxyu6zkb6V43L/Lt4tLZAXShzASUkyCKKlJ4pmHlFoYtE1LxehB
A3g/aQ+QKhwO6BBzdi/69apdxC2z9uSWQiiVPzixaLqkAbBIbQS2T4D8dMJvglDhoyPxyXtDJfJj
y5/nlzoSM8rQD3whKz3/AuhrB/qaUI6kMVwIbhGdPiYzL5fMiEsxGG7N3PT3KjVlW/a/+TvzuTe6
46WrGTRw0rwHcWCfoTOf0X3RlqhFn1CMRr1hyWam71Gx1AUOoQxVkZ6VaXxa9dbebQvOY4PTrkEy
prWj9JY4tlNaEWSzYaZWqNbG2gFjvHEeN/2FJsNJV7mrhwvomkye5nG87p+lq+vTTNBoWG8Zkkfl
unV4WdgtSBWE1zAdThqKqpicVXvbWZejnn266DNXZPyq47iG7qxTBKf4TqoOs1QouI42dWBr/o0/
IXxXRKN9n5nPMK8QaEvq9qrCeUDhL9a7W1RjxebRChCvBq+Mf8WeWzuqr1UeChvYS1VuQuIPGdRo
BlpCLRzeL6ohflJeHfhZcMMqC86Dry8hW2nDI5FfuoqReueshgu+ufKf3voY0YTsVI9E72BeJtuH
rjd9dVR7OdGGxvfMEAPc4D6nB+fYR5z0Py/NW/l+ZL5qri5pyPyYnSBbD4I7Qj8ACupjbimdoPf7
0tDfyEVPOTotAASxInEJl+PtuuvvzKSb8BHNcM4FRH0rmzhJ6FicQIL7TF1EK3ZseXZrU6LZ4wod
+zpJ9PAiDAc68RjgiJ5BDxv0mmu41cMTXNjWbwyFzXRQOxdkGdU9W/yvHbJhXsg8qNTX7IFnlKsm
vTUVJ9vcaw8inR/aJukLoapRuqgQZAP1a+34J6f4DKEjkMncuxMBMVdPKZIVzCj0svgbCZSypwnF
VK2PAOPj4qDEepdoiU1AGb1dgqURleLwt1hVp5SZns9GFCvY66c5/0HZr2hrFTQWotKggT61JJgu
JKtd+205TTTObu8L5e+3RDldSlJLvUSuE42cuqtLkS8WG4DE4xShE2vBi0NybapRo8dRty7nrPpI
8cNMmPAZyX3fTTAYQLLptHp0KPNQ8eXNJlEuM+ue5VoxtxCDAnO/lcf+2aplQv//oWDtvhpX+L9q
WQDRKJe+M9JIeM0iRRHKILveym6nuWemZQfqUR+eOmoGqxDf+UtnMTCyAgWJLHvmyCq4aY2DzwI0
TCihMicjG/3oA70pkfbjdZfeK4ayvu4ZGRs+FFzdTZtDX6MPIbhy41kdXymhpoupfJPLCf1YlgpP
kJGmMHqeA5MocqKLN7SCUsPhDhyo1j8KLjU7+E5pKw9MChXeAO/yclMfAzCN1BYfEbf0tuUmJYQo
Ou3mXm0CdN3freqfLFQRB0FNnnp2P1B52Y6eEn+Mz1BIgUp771V+sbijwp9WHbddZBuEfQHvBk5m
IZ+TZyxOvg1qKQuqJiDgdGzmcr8sNt3SFNLdXFTlhSozB9uGxD2ROCAbVRLk+wHDb97YkIjSvU43
4ne6GYCP+b/pzrNE/ZC8fl3lJCi313E1h2yBRoJNBn1uQyonQGWc261Prrv9dDxwMR8zjPNbLoQp
FBMWvpDmbZrKa5Lbe8xwJZOpxpcZ+bBfjFWWi1VRjY2p0bNERQvnDgSy4RBCV1kxuQGX92BsRLzN
Cbbb48raL8oqkCyrmPKb58QXtJOy+zrImov6wUOvudIAdCCxC0BWnqelkccATa5LFGQOu87FTlQ3
GdvLgkT2aK7t+fIiDnTEUwkkjh56LLseSqr/bgZQr5AeGDKLaw4YPDlaUP0899i0LEiLcetuvToH
gB4GfUIW4v6HEPFyVq5DijYaHLggwS34S34TbH8AtTnUkZf/TBzgxTM393lAauNQufn/M4yma26z
LoA3T3kq5BSCuwvnbGojV9ZK6Qs9rRV8MoAUDTPU+vL2GR62Vsf9UtowtLF9BMswLq8BWBTZnokY
dF3SFGn4+GoOmg5LLlHyrf/fDq7NDcFjO1/r0X5zEhXq9/nhoteuNxLu17mWifinA6h2Qfl/bua1
lXrablfXE69oiHa/6cWVyD4DaKv2RXryYykQR9DT4K9BRDj6yNzy/k8IBqQgxBmbl7MOPHXvHptp
hzKraHoCn65/mWkTcPxH/k421TKCkG8YL4OdArYBox2Av7ypdxgI63d6KFhENl8ZTS1mET+ksv+B
RWMWDHpZF8lZjGiN6o4m3SdxG+D+O4onYkFd+oeRi42hHdx6t2JeqfuPnGGKxkmtePWvuaVDPU58
eHklj5BdehpaC92RvFsTS/6KL0VPIGBETWM8Br6OdehOnXf4Gh+RW8pN2NPRhfdwAM03jErBTZKA
+Qpsu8TFVtodIwob1Wm56D1bqOCrR3QpVsVDg/P/TSUAuVkajIbrOVeYYiCVNEpnrKma2SUh0hsy
fCL/j6NXMh3+e7aNcqFXq75g3r2D9uztnoLYw0AMJKapMJglfzlacOhpInZe6/VFmj5hL9JhY8CG
Wc3RZ+p9q9QRZyfSrOOm5r+h/7LEgoswfJy096hBmnXykV63lfocDZOkf4ooAsZX7g2T00MW94xj
CzYAPP9/+5RwsIQPqbQVXcpA6pxiqdAQ24KVrUZvzLLKpF1wsleyHrWxDAmEbYR0dYTS0YPnjdQ6
2Tr+3t9vCfLZKl2asPwGA5jTbkzksdVtWEUE3A1jgsdt1CFJ84bd7qOrmgJKGmoWgmEivnHBlD5t
q/rS7gTRD3W5N/QfiSompCECUiXwUBOWQThe5Y5BVu73x74KmXjKAhiiXn51xm/hKkJnhgrArafS
s3YskHPzV4dy3uASi88g/MvONdqSo50jrZ4Rj9wjD/XwTLAI4XY+i9Juwszz0E7qxf5Y9yUFfkCk
eGaKqOtBr6amosBxp6EJ9sCS74rv3S/WWJdrl+vh5eAtRA7DwwrUVlIwy2QKjw+AWOAgAliE/Cw+
eLbMxBb8N7NePyo8SlY9vet/U71xblVmUbdt7bUmTLsL6lnG1AOEabbVdSKcKKt61HpQ9+ynBX4A
ZMbr5k9neDXXNINEF0AMeDKfrRkBd0MrESm/MgAFmKsMRcBZrS+EQyRr+hwVDmRrnzj0D+e+IXQ1
uXtErQZJXWqvTCOM0Xwfo6XMJFsQG3Wv9OrZBrHIwhRxDInsz/03m22wquMzdw9vlaYtgfxa2zVt
S4O+YLgpmu5TWVImotZ9qqunequFPpStYQCIPAtwp23zleiqY+NOETcvNg4S+y4yrUCMvKk4jU94
jvHclaXJT8rR3LRMW2GXiIp6x0cUlPpJJbona4D2g/9uTUdl+rcPA9yJuuSlZ53JDAXgOa28hhOH
hzmhVV3MmR0Vx1QELUg5bvxMeAXN5dGvFWBCnOHTKHxajTZRmJ2b6a+UBX1BgSp9+e6JY8Ne1U2N
GS0wrJVq35Qv6RmMFX802+waQrIEmO+oIz3olPA5pDFJ2eh51QBkxAoEuEMSI06c8NVUUkkSSFO3
b9wV9rtdlWvEYBli/FfPw1G5M1Kv5gqHNMZdAuZNzvdTvLBIpZLlj+U6Idw4KGq3GdRnh1dada2y
RY7WMchme7g68M1k3JBueMi9+4B37f5esvIxtCYEQfVowmlD/aQXYSwVw1XYxk1/8OefBFIlsNk/
6k3z771EAu3yPd30KdVBVL0f2QFCVOoh/bUE3fPop6Sxes9vSQEs73g80SohGYykWotb86PyutKC
qDhzVQQPU0trPcRp3T89MRL8TRdooWlsWz64nWZcFePaBxpDhxLG0z+7cQajUZnoOVFuCf2mnJqv
cyuTKVKnpNyV50rz2Kj+BCFInkR/VyujDPJ/xkD1q0pdNbtqy9H4HDRBzr7VGf8UC2I7tjtWLeKL
op38p9P1g0DJ0szZWwMfdRLEAczO3jXpD7NOU8poVp88ogz/FPXq28oeDp+Ak80W1XVYmefqYOxG
VXPwt5rIgmoC6j0GSDMYn1bfytcVwtNiQINKFWnSn0qWKkSxqzp6R1oBZsdC6YTLmotEz5D1dfNG
6rWTvkchCALp7ET3or63ejNDcQHHF146LUgMzF+N+iLSRYNN0eNnmHed7NRf+lcpDrIcYRLT4Ygh
ZVfRgVK1JUYiWdSHmRHT6Sqqx7Je/RiC3eADNRkzWWfn8V8B+YBW6aLdANAHYY2Yl9cQcbOIpZez
77B8kN3Sm/7zlSbbg7BZgPUDwEg7OnJgsF1r9OSwmvcymnolnaOOcGGGxGFd4YE1Kul/OuaMPNCo
N86oeEbUBdMuK550s2HWeAULRl8zWP3tWEV5kGA4BegakxCu9KAvWBkECghU0jD/fYu/Co2mhQDo
z45fT2S2ndFlfYir5VMZ1Gn9VHK9CxEsP4hzy9No9X9tjrVh2+mbfWBvYJvJ5n1RwSco9j8LZJrx
f179xv6vDJlXYMrQ/PXCpHWYwnTFE98TjMDO5DV9WAeoyuJLEOEVv30KBaKTYmxY4OjZ3wCRRB2k
n72UwCxSXrlU9Gze1GaIOrBH3ZkZFDdKH6KfowjB50TGvKZtiGTdXRBnRzNA3zWr3lxEoXsxfuKq
gmQuADhSeoPv+P647BRTnHAdUVKxGw6S5MNRnUtqloYBZAKsImjyd1MktYzxmUoOyYOsuNBcqSfi
L4q1f9Rw43n1xB8VOe17kPGVkswoiyqlTCcV7N8ZKN7JuAr0oxnX5BUeeApIz9JU5qy6ZtzwG9Ko
7nE8GkJv85Mhw2TqqZgf8ZDI7NdPr5qUgi8ZctpgndS4r2pQypJdibzwjjjAc5ifZ+LPTAKEyUPy
xxa/Se2fBMLmXqU+A3imVbmP/vLQqXAjFaz2Ag81p8B4J99ElQJXwIWsYAiVn+bBe3h6TypvFNPO
SemkrBzPMaOfC05oz3gKYVFsD0OOOrF3g4Kcb3cMgS7Ll0m4AKC76HPVM7oNjapT3CQ2lVLA0nd7
UrdxtUDRUhR+x03jzkap/E78Wk2H6n2xmAs+rSbH6sx27JUvPVome1CF+YXLT3X9P2csIoGmlkg+
T29oVm/oWjs2jkcuQC/QEt6VAaN2wRps3TPhtMwu/hAo4zusht8f17XVv93UvoiQTn+6L69E5iHe
5HiYPwKbWMof8jyxHp5aCksx4K7w1B6kkpEodJ6zKuw41UbVNYYRVDbuPgJeO9h4EzDhZswTz8ds
eKwVZ7ooRlJw6VZm2p9cc+hQPSn9A/MGSAfKoU0BMr/puuZusH5CreeUwO+4btHz5SfcJCiIhgl8
SDjsa8RvPf2Ce+AQ1SWTpVrxKUWJNG1/OWy3xvUd050Zci05JsamKhFVkkImPs2NllaLZJbGP+/v
wdOJIa+GNnOTVNfV3EokWrnW4hKNha+F5uJ0HbhWqWVE8ay6KEeGaPdSgp9GjsyQnAieN/AbdaiB
vafPuygB0nZ7ffACpsYawBYHx2fahXXxszfpgUbvPQgUzRNz5CCEIGRlzvBtr7OwvfhVkua8/CLA
aByqIxYU2XhtAFGGWAcMmu8mrwY7/0ZlDwvI34CwfsCrEptkHNSsS7TEZAV7LEQ1McZ8KJ2sQYTT
tT4nx+rVA2xHzLRgEBLUWkDRucQd16o2JNlGeH1dzM9PDQf6BnbGqQgywoAO+O+50qn0y+q/067p
XQmQQmlq9e8SC7NqqNkK+OcnmbRnYaD/7XskwrYioCqYMg60qeTa6/FH9hsn+NGRD6JTnFpZjAy5
0e+8lgpRq5OguwQaJGDLQ8uuhksWdngT97Auba0DsGvwTQ+B5DXr6xxebup+UejEx48tW/SALq2w
g9OPzj8I14NvvIe43KxZHvaur/+K+3+5zaGsRcAvcx0tultVTFGmgFuYflC/92NzEMpQLn3yF+ps
JeljLc2uiGU38WgPD5qV1Up39/FQE//ss9e+h/0hCncCQkaLyC5VcPXL/J6aH6z8kuY64NL0npQx
5rywkDZ19YtoI5aeU9VVbF2rvX3wczD/2kIzHZyIt5C7FMVnYMU5Rn9Jnnc39VWLve4wsmKEAeRK
0kVV+GbuZxzJGCq56xt5Jq2eOgzIDmSwX5IXYMOTabo8CZJuAigP18I9LE7coq+iWyKIkA/2osoH
GhhrtcDAUWUfBMX2pyFVgPvFOlIpQw6F9hKArQsoXZsOTXzYmzB3FNLpupf0SRCCFmOD2NSWXVo8
Tn7uZO0A2Tap3+CauRo2wu96KXZxfnpjiGXaGpXjjVCf+bTSLdOE3SJ45RVXaHjJVfUtq0GLMjKd
J0Is2+rdAT3/er27/TJYT20+ThnjNtQ3wt83YT+bNSOfUhQar3yIB0CDrDu9BmgTWXmYDXW2h8MD
5d7ouVIjzJPT6mz12vuyorth/MLITYRVlT1DcA5Dkl/xtrotveuv6/2C7B6+gfQaIWpFHMkJvk+T
tKkX+mAoqSbjvt+MHp4V0p6RSAjq28jy07vF56wDMNUPAieeQctj4XgIJBQEKh8mIlvfamTui5wx
LyLvYzPCQVnKt2FOu9qpiDFkMHP7KOGaxMxxPJNhkWmCl+OgkaNoBjwIPBoFb0OXGmqwl/FK1TVR
a8VZlEnHBMVuNj+j2JIS8/S4Rc4ubS0oLdVIjXODgOJVw8W92giPzju3a4IzWrZEtxytcQbQjkVT
DqDpf1ZWGpIm3uPr15qrTD+OEfO6XSNKoJQvBWbc1Ab0dKpVD6IKoLCac6nrWwb1SybvejMJiRQ/
OJfr/1jl/lui5VsS1JMUI9LVP0rq/AxzbkMKnEAGEgIIsXm0uqvtNsUtbMHVN44+FVfDDDf/yxPw
Ky3cv0szk0OJFtRdYaaoZO+gWYemimvpNizKQpc+q6LuPPhKVH5MYGMHVUbVFW08At/nhSPr7o8H
RmzNsIt3tq9w09iqYqF5FUcxlgIGxLxK9j4UIN8A9riXwlPWmEk4I7xAtFkCxTMyWuxfq3CcJzHj
MYz14rNnmNfpy29bHUpqJcVUjKLOUof3RkczzNSFSWNwtD9+iJkkWXPF0YNtqkK3e0l8I6ypXxJ3
LI6Cvjjs/EqEBbiQA2lMTL55vku+MfNDI7ZJisek0PPvP4K6R+QiYRD88vXSU9g9lZ3U+hGn1Wls
NMLWWoEczwUCae4sz2mPMSsKQUt90sGEIVcxRCCycaAk6gYj6CG9QaQrNq6EcG+oZRfdC/hJq2Rv
U551XY4T9TFPXGuI/ah2QrlOx+xUMAUg+Vs2qMbMw8d6Z8Gufxqw7ouR3dplafaGydny1U/Jt5OG
By3HaR6WJc+/xYksJbg15O0MKJIjmbkyIFvr51tO/EECohhtkO6WGHFnaJVZ1wJ3rQKsT0W7LwGC
cXuMk2qJourdmG7y7Vw0ySoxCvCFvxn1ExjTzXtuzHCQPHmt7zbdg9WpDEROIbkJ9JxiXeQDOtax
IWbZjyuF5MC1MRpTuCgESSMN0rjHWcdoi0km29/uUh8bYUHdYJVjGc9YnE2e2dNd6T9L/7f31s9J
8KfRfcP36ytRzu5aWahFTdRMhWUtOPp+9FdJVFe7GeLhj5bo5oenrAhOyKPpdVl5K7DTK6lcFWfc
FXLACubYc0YFpDbVPFKMq3lXzoLEqNK4OzsnkvF/SgzuJhSujeXojrbDBSpDf+xu48sxC0Bkkgvv
Xhw4JzYZcjiMVm73uNpPrtKJzhnXfPw4yMQTzKFNK7ZIN8pInjpL5/sueN1j03SdFfudq6bKbcv5
oAbKK32U0p6hdhXOlihtzZBAh7aXCga7nQnTAH3tadsIyOHll+xk3Gyf1nrjBCxXJf1uTOhtUDv4
mLS7PEWdJAL+9LlpoFGPKyzhGfXyLgmtAlVhEoO7WOmkEjpD5pnJirFGL0W8ypz4a0uQ6ZbLniXy
fiLUOPpE65lqoijnkAMo/60nJc+VXvYlQYM6RKLvDl2sWAd3RaHwyezRU7lmOCND+Qh0rkB4FVYO
TremN6YMQydJY3JBwAtOA1FfOIY7IrL8zzYhM6NlUdp5rDXDqCwnuKLfbAo7Z5O6OjWqa6O/BnO0
GCL2Za186/gXyaOmTEXDbqwy3DHB6h3wvWyu0P2QQkmsK+6o1TlTxp53O7NPO5heq3HpegMU+/nv
UIKfwSuKDtC/mGi3/EjANEfpIJisz35ZZPRHtvftMUG67cz8xRey0gO+ivKV2FLLczD0VdkW3BQ+
JngLADkj2oK1+O4W0Xy6S8xq8Ok4OaF1VGobdiTk7RIu2kGOHQPCkuozbTBU4tO35jzuuA8khD6m
BPFXYbGW6QvwoBcKn1n97x5sHI+ePZ13hmYsoYTCoRMs161ESUYr8UD3nfCKDm5YqRUOJO3KRada
J31H5Lr4Jt8x4NExSSU/ghgWsVNZnN1QUAqSshddolQKtZXk8C46yLdbWV0KqcJzrxp+yeVZvdbE
wgPi6yOVCjxTRFWNzf0zaXyWMD/u8F+fwrxfkw0bj6Z3J47mx8kEy5vnZ2UGAInwKc40omxlQPQo
sHtEfmi0LhTzJF2ncWRQ7Bm2GTUzXGo5JnUehka030B2AVdVb97pU2lDvqMa5RqJBU2KVmbyZLpw
zhrEs0RIlPkf69P5sIqDtvjri310tF9pxOkrQbS6OCQpx78HQzyFKjBK9Y6RsZ0uRnmkFI1vDdAI
vwMHIqQt6g0LIJSLjUiB4mvI26sJJF/kzIzRGL28u7WXQjAB+K+7ICpVt8t/pWhwnvv10/fleGBy
t3Z/59fu0/NDpWOshZ70T8vtwslSE0BEjr0eRbW1rAXUPflzUbduPdTAmtxw7hkWCMo62qoqkm6W
jnRXPucLPmJ59qaFfQBu6uQ6ipCiwYA2kSbAsQ+M7ucvusk4A4SsHgQKW2CxkppVtwW5yWKDg7ke
/j0ingBnhPWjWqFYKQ23JDAc906rI4jsm9GfePIZ2QjFb40p2ZDk0byfYezzxrZ5TDdvOV6xt/HN
OADPnEmJ6cAPQ8lcU+1UR9/II4crPBjUJ8rDJdA3jsOE5xIg3GQNWGa6eFJjsetDkMQqo4kvU6Z9
wNAly8NVMIHrQaHbu2Di1NITZNbB5rA8sGufnwQ2qDsv10vRXmWyiNCti9wtMMjFCicK7i60WT2R
4Y+K/XhPRxZ1SmndgT3nXvnY8/BXY782t8U7kIlmdcqbZpHnjJzkQs38gVmKEYx6nAStV2ZEzdd6
SO+RESSLVrdp1EDpfkiyiNBdiyURemFtdGRhWENfaF2GKcPN43mKQKzN5HlmcbDNkcvBOoyQSnFd
ONoDMYnVEVzDyxyTHv9O7xQxjN8+vRVoNnJc+VxUyaBDHYVGfWD8AD2uyUeigezcebVbd+PlH9mS
yysy6MVZzD9a74DPcOBKeAL6Oq8xAIgR2fTf5VGxYz7aJezLSNCVt6zWsPitAektf0auH/S1QFV/
PRjCJtZBCTAnrywN271R07PyUpzoViuc6lmlqYo1w+LUknOYdz3cGMf7+thDF+WT8cxPN3/aKNNh
Vohbx/AVzIUb4XQoG4593YZfYbOr8+7dLmb1CV350EqXzf3YybNf3d8jELw4qxGzOf1dUwnZd8zF
XF1kmLj5vRS2qqdBKgDrLjeJNwVo9JfnrifEI6oAQDa4RSm6e7rj3tAx88qYvdTCGWfTsjLmDjXz
UPXXA0/vkl602s/75WYsOoMwZwRnWHMpP1vjOj3TqGZsHlECoHar2jJGIyvZcgJi8lfym+vthueJ
qFFEnmrak2qXLaP9Je6NNqYoaRCBGvrNYlaJBW1vlKZhHpO2i23a2QMrgpXdno33V80Ngh4mEvrj
0HViLRpqDDvx/AAYzDZEsLYPwRzKFiMTwgYi89jh5ML8fwRaM7PAcpCa8F7YP3DRxq020s2yqr2j
aKwBPhQmMjoEC/jySNheCIYHNYF0M7TnNe+nNN59ICbdX0Af+NoZaPmbhBmj2Ltvpkf8UZHXeRUp
kb0Ft6s/RWXK3SN4YhdVtcXrCIDct41h1vUDNby7R5pr3sHrPEp/yUWkl5CQDr//Q7KWgUf8db44
IL+XenglxJ+xheUFbuqsSiQTVekGjndNggh6vAXj1N08Llq9gih8UNFoeiDKkMLnxiiMwe9rtfqs
R++LOfxs/BQctY+LahP+1gUpZ2BzcEok/4VY4o0zcKzjwUQq85L0CI3mqSeiWQ8zuFEA5WhXFYRb
HYkBpm3NyYnlU7001YaklL/TVfVK0QsoPhttLtyfMdxJ43EXmvpoXQj4dI43rEOdzjFdm5/H2jEU
mHrc3hqLbGa0guaTCz3v/bT4XJbliOkskc2glZ9Wyq+L74UV0Mfzejrtu2xgTEyC6yeehpW7kgzR
ZiTlprbwSLQMd8ttE5Pcq2nPwm1KyC4LmGJvx1C6kWC7IfYUn+JJOJ/iFXW1MNciN37kFRs8F6Vg
dgHbPOeHXablm54q8nEU+5hCHYK0arQs3lntjh/lIJMx441ZzDMu4UsffukW34tQovvsUZrP/XCo
IzIDG2v1yrDJJ41YhwXUp3FxhLZgzSVS46QyWOtjMoKvb9KuT1UDF/cmsFI3mbc4E1gVL6a3SB+l
7opzq+l04G0STC1ve7r5g4qgIq4C54NvPbekcB/cSmKfb4IOcLDac7O2NJCBKjLGapHn9OXi22sA
bQvsvm0TJu52ZECTpYExH1KV1ao+HZaW9o2hIblDgu+fWj8XImfj0h1CTPIdPLc/m8rKD1ICi1WZ
K/AvxqVq/KjhCFYzw+Xz+bj4WhftfPKjAdaZJZFNmhtceqslGGVvnp8Ya9/00xpNaQleNgxNzc5h
K4ZhmKDmiZlXZO6GqlDv1+aooV9qm0Rm6WxBSU3AhrJJp6EsSGmv9pLh/38nRFMqtUTivl2XEOWJ
KSwlHsvFn6ubpS6dCqphmOjjtmOLKQK/SNATs1VhD0P/kO1ldnPscyqeGOm+XR5lUT4vvO6r/76I
kfpy2PCVGYK3o4ZwpInRXdYxBe3McjYeZNN0k0lJU/8kdTn8XeD3D7M1eum7ep0gxKb1YLyJ31bJ
3p7iYUeMLj5bZQA5sZ+jXcbnhQd5WUEzbQIx/oZhekwtjXngj4WXbdRnXUv9rKJh5qLrji/uPh5n
ZwUTpHjQmlyGYQGYrgPuKHcd4nAAxoaEjTQDFKzYKoSyoZKXf0jqVSVDv4/bE80t4tvfdm51X5we
56mQvVyXKvupd7zNONKKqXKqm32lo2WI6k7DWh9mymv2u/9yH26334aUPeLV7/0yba8fLtfsaq4C
EU2Q2wBvKr3/fyEB89dhWu/cYt0Y7d+kDxlV7eWat5cie5Ya2323OD8JxgsjPqu+ZiYNP0jUEq/6
epDPhGwdKdOSBue45e/9NhKxoKdxZLGdJitMvGdFxjTzJv3Ju48MdhwxvuTNI1OwJtUzE9RlEzv3
ucD8ywOLBjgWdYghXJatVZPTwByQ5H6s6KDQVCi8U6fJURnVrI9ZRbuwTAlV3AgREkbuhdLDv7Mx
+ooh3RO9lYpbR3fhyrkg4ysg0bHTuZv42byiH0Oh+JvupFZO/RukNZaPc29/18ACigVDvqyi1wOF
J9at+0oVcOqX0qHOO63k1jjLbQuYalndMNwHcbPCaZ70DQG8ts6UrW2hSqwKzA+F7maZ5jgbHH+J
tGVoUQFwJriISeMxo5KWqtV6jqrzufYu0BFAe4oPDw8kEaUZWqnvTsCDvZsDyYHRmir1zynZT9I8
7h3PkbDJ8mb883tLWa6tD6IhlZRnvJnzEkY//rv8Az7kd17y2dpXPiim5U2cllA1xrSNqRExc9ud
kEjm2nZoR+bjSrZESg9mIAD48D/mDUaX
`protect end_protected
